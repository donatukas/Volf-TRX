
module DEBUG (
	probe);	

	input	[31:0]	probe;
endmodule
