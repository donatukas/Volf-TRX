��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.yu�=�6I�.�u��)?��"a~�w�ӌхu<c��4�<�u��h������=`�y	��bP_�MC��<��\>v�$m�k�q> eY��N��n�]����`9S����97�c�p��J�q� ��uċX��"�O���^?\ij�7Ƹ;(�a�o�q5}kфZ��ϭț
[���<��w$G�[�zY��g-��cz�Iͱ0���.oZ����\��.f��K��ש���~���L��f�oO��u���\v���]�K�a�3epu�4P�����uJ��G����������.�K��1N�X-R��UF�T�䂴>b���
�'#~EehL�����h|�v�s���ZY:�#2;}���ݷ4�x���y-���P���c��)r5�;�{
�aNqx<Z2S�a�؃�Ć?Mz��2/���ϋ����:""	�p�d�gƁ?K@WÆ�x�p��:ǂ�����|���vM�*��ͯ���`ro��#!'��W��e���w��;���.�7O@=�O�B��c6��W>��-��抡�A�$T{�R�
����-&m�}O
�����7=K�?*\�p\I�{��0,�)����j����`���X l�mL�+U;Q��¢�)���^�g�}/�>��f��HE��C]������b Kj>c$�RA��+	6	GLit�	��}���Y�g�f��6<��T�Z&��E�ZU�fl�,|��JΏ�e���+�J�~�|����390r{U"1�w��T��̌�ɕx^	3WMz�����^��O[R���'c�*�.�_��q��)q��m�#���pZdc��N$B�U�c����1��+�c��C�l�*6aAE1�����̘Sˋ7Xw|���(��R�����=йLǌ�b�|+x���%Y�y�0ųT�����<����ePG��lDx��r�6O0�����׶�������ۣ�8ny����?�&&��Q�Ay��Z&""�y�v���#$������� b�od|�&q��C���f�V�!l�ދ�.FRҗ�D8���ՎG�`=
%�$�ĥ��XP�/�������0C��z���wM+�n�>��$���*�Vt��&���v=�����3�3�GCC�t!�֛���T�!�wU#�HWW��p�=�0���!�Q��G&'%����LYJ����
%qv��lL�k���'�Ayl"�of�FS�r}9��f�\�v̈��g@@ ��x���q$�o�N�T�2f�jF���=��\�����Fh��6�������<Փ��<桎����o�×���Pn;-����K��z��W��ܽ���DK�3�$# �Rk���!���X'�>�W��K�!��
Nq��'{��]��	Lhq�$����̟�2x ��5-�h��}�Y�ģ�5"���m�
q��+?��ܤ]s��ƏO�K-KD9Y�i`�eQS��y��yYo�	�$H�p=�R!�>hˈU٢����a5����HH��)G�M�`�MYC�_v�-]V#oӲ�*�'4��ُrƛ->W"!������=n����W��+��$��Ϭ��@�{c�
���@?"�ޏ�f�"��a�dK}w{*��H�C�l����8 ����K__�$�xk�q�H���4I!�
^@������HS4�m��[��YZ�4�ЧEPbo����jȂA�v@<��DSYN���9�/�Α��O�άeF���_�h��L��QB�aԾ^�p�UR̞����h��֟-(|i$���j	��븲�#ن@ma%i��5: %����o���w�nM1brM�J�5���p�>�?���m5���o����[�Gݖ�$܄>[Rj�rxL�c���A�Tes�Y�(q�s�<�BjsA�)ty@L��׾� :0�3�a9�O�{5��\7����)��w?O�� ʖ�	���0���Q��8x�2�� ��� j�%�ƻƀ�?x�w�a�M�
Q7`Y	K:�n	��$�g~m]'p���:Q��h�C#�����Kq��ug>��|~5�=�fl�������R��ڛ�)�-+.�n����$[Z�:l�]=�&��@@�D��顾��.�c� �;���O `�ch��$��1�is1�T����.peP�|+�r�֘33���Ƣl	+P��r�4�u�1k���t�"Y󲓄a5�R�.�~XfA	N*=�l��a��Ksa��{52��/C}����%^�L������~tsH����#�y
��T���p�-�#��H��De4�/�,]Qbl	͆����ۑB��h�`���v#Wgy�Y�4f�PrmH��;�}hd"%��|�ܒ���NF7U#ph%����`�i]r�f���F�5ڍ� �C��
h��������Kֽ
�L!��D����\��w�r�P;����Wa ��\����k�~�&~��[�+iЋ설I�fDq��i� B��6Dx��?C��\m�Ϊ��m�p�G�eFW��K�kS���U)ga÷�G������R��p}�P������菛��9�
�����f	��irF�Z2a�`D4�:/S��UE���g"ȘJ������s��*ۄ!��]�\ts�r8]�3��kF�5[�����ץ�a��yBr��8�뽚 ���*q�&�,3"���#/1���ǿ��,y�$%)�(��V���J�o�(��曤�*z�x���̽�)�8�F���mi���ȃ� -w����J�:4OdE��7��Ų����bѵb�7�+YH���� ��I��&=̊�OsͳI��1�g��b�hN���=a��屿��S^��n����l����X��9�p���N�kt��)B;����0 3�6㶍?}Zme�y,$yq͆ۅ�����8&-t��sM���ܷ��v1zPN5Ƶ��wn=�a3�u�I[���#�<"P�GP
����L�`����Rw��@�X��6�Aoa�Xl,�Ǧ!Yfϑ���t��o'&g޽�ĪZ�D�7�K;f��U�^�Q�/�WZ�?�؛=�����%�����J�:y=�L))�6���r�w*~	#��k��プ�	����儿� ����9V�@z1J��4����59+���v�bw�<yg�{��c�{�ر�P��R�k#ڣ��_��N1�3	k7~n\��vh������]QɭȊCЦT�F㒥��]N�ZNd����C���hjw�����#��6��J��~71Et�����"���+i�M6jq^Γ*/L#�ե���p���V���9�����D�2���T��/��j��r>L׍�����x�+���f�nJeT��㮃�e��2dX˓�`�+����Ґȸ�E3C3�?�m�T���9p�]v�ϟ4Nw0&�D�8&µ;G�\L]�g�"�B*L��0tz��,5�9L���֙�8T�Rl"Y-b�j/���x�<+]m�Ah݆���2o�O�ZP�7��΃Iw3)n䳝�7���9%�o��o�7��#I���B>��$T8�w/�^�9s*ܩO�#T���.��8�[���&����'��4k��>]ݛ�E#A}�@'��̈���olg�>ӹ����\˜g��g��j��EфS�5 9~三�/����@Y���^�O/�i,�:3�է%i���UB���2������D�w�q5�	���1/�F���;��{_�m��+��=�r��ּ���	�ddc�L�5x��r�CS��Ӝ7wfj�<圂:�z�g?KR����ŀ>�f:��j�M��A/0jT���3���:�!}�MlD.^B�5$�.��"G�u���M!�i�TM�A�C��f�ȹ��n�'�2@Nh�[�O@d�v��	k�z�&��T��s��8�*�(�*�x�FQ�25�zܑ�r��H<r���� %E<�i� b����������4I�����~V���`COQ�ӯ�!�8C�J8 f�N���P�����.��BW[)|~t���$���ͪ� ��Ml�-l�ta�ݬ�/E�n�>X�sd� NH�8:�ɹe�����DrT}�C��p,ds㉅J���f7F��k���Ⲷ��3[��I<N��k׈1������p)Ɩ��$x��������@� ����C����1_8	�L���g����Ug~�9Ă���W��̔��-4~��gˆ����&���Z,��/�Xiu�4�J���H�ZAp
�˚S9����H?K>x��
E���4m�=}�v��[B���k�v��x;lD`�r� kXd����2�)�P��P�G�E�gT:�3���y��@�"
���}����K��OU�6�{��"�u(�Ќ��fiv `�fbԯ�]޳X-h�����H�$��[C�:��8�����V@�������P`-o�
�������o1��|6���D�9�#��@��o�s�~��ai��]\Z����C=+
G�Y��s�D������C6d�Lp2�6S��ǌc�x�yc�>[�LWvZ��J�1H4 %�r�z����R�Ir �R��:iu���>�OS]���}����y/һ���p�:I}*C��wO��g�#�(^r@��*��ӹb���#[�Y��b�B\~���#f���	��Qk�m�쑀nB�Y>s��s�J��� �d��u失R47G���Y�Y�n͵I���hp;��T��*r+���	��';{�<����(�yg�;����i�XH�@�)�ݷ��?�!6�5\iH��y�8�8�h5�#��4��&#�u]�{!�D�͞��a�3�k~�>9�+����-��I��\e�͠s)۶^�{j3�^2��CmA�����1���P��ˁ2u�5��q�&�i�Q��K��z��="WS<�,�NbcE"T�������ޚw�hu���O����<��:�����8����7�F�aC�|���%�T��Gd�4Ǥ�l�q|q��?�X����u��F�"i��=m����s?&_��eZ���>Ab��.B�u6�2���&`�ǭ\CJw���s��\����&�<��)�"hG�*)�R�����T��� ���W4��;ǜ�h�9Z�0���HW`�'x�5q�h�H�K�-x�u�X�������c'��e=q��i��h�h�i�Δ-�����`�E<)u�l**#��6&{e��� ��OU+�-Ѻ8�8�{؞A?�4��P�8���˜��V���$�l,-��߀Z�pS!�tc��{�@(�\�������9���=�&~\�y�-��VI"H�'�d���l&�0�zTߦ�2 �;n=�-��V����x?Ci|��#U�>r����$�����{���oZNID︕��������g�[�Q(?'f"�t��!ضď��RєY����zmxL%	�.��*8���[X��؂�M~5�ir��Jy/;ܷ���/���-xci!{;��d�\,�V���hZ)<���ߛ��gUw���	9�e�3��`!-�X�.��Ro������Y��[�ۊ�n�Y� �H5��D`Yq�K�=�P�}:����Ȕ��.��6����GG�l�^�ˡ�n^��֛'�~$;������`&�?�}��\od7�l�g7]E�$7�TB%����b��#we�5V"����Lk�,����g+��`�1�	]h�(M����ģ˕�B�g�U�Y��K��f)�F-��^V\�H5IT�ζxuҖ�kc����䑫6>�tBJw��gZ2%�r�|?:��P��ca�<�O0-\�RLv�B�x.5�Vž�-W�A�U!w�І�xA���9\���ʺ�6�������Y�-]U+aU�|Vw��O�:Z��8�.- 	�� �r�"r�*����RW85�p���3~ña����Ua�*���q����R�7Z᥏4�\C�'*y=�������n�ȽN�")�W��UgR~� �0K4�>w�v��(N@٧Nn�{�.ƶ�J�+����#�<���E�!�"=�/�¾U>\�v�uw6�9�����m�l�>���W��S��1�u��9��:*f*D���C�F�cBG.?��MlM��6�
L��y���M\�W�	C��8�>b�!�?���y�쥒�ʃ��@��d��l�ނ
4SWb�B70�	�g�Q��/��R�i"��{��f0'������xMkF��e� l��o~�Ʒ6�u2_!���ڒ����y�"8�j�B/�e˚��a9T2��@a�[�2�H��G}<:�Oe?�^|����n�3�NF��\ �_P'ڛ~F��S���h<��3��A���R��X=,�G����S��@O���c���Y�6i�f�� �w���j�~��,F<�h��D�|�,��D�CԳ}��S"O��2,�K&sA���t�N�Rq�@{mWn���W&�<�5]�t��]+���Y���"�F�V��& ��c�����iZ|I��\���?s��n��L9<�DșJ)�}�ܧ^EL7;آO���cx��!��Ώ���ݫ�')&��ê=�O��>)1!4��Y����
j��x8?.���Wzh�CpT�o1<�Ҧ��%�������kT)	���v�qw˝躝�ʳƙxNƹ���ڠ߼�L$�Vߐ
�m��(B��o���L�Ϣ�W��/N�"��'���J���;��6��WЫ��%$���/�y��+�u�bZ��tK�6�F��Fn"�(�w���DO�턛I�E�̄;��m�6�:q�P��%>��yBE�O܀(�f$ļ$-��4P#�mADu��-r2]?�"��x_��rh ����G��	�����Ｆ<�m�ʛ�����fV}@x�����i{J��w\�|�i���a$ s�y�Q�}�LV�f{���_��w�g��G=޿�o#���ү��{.ͫ�O��	����"���y<~���]�P��T����y_0����J�3�<W`�/S[�|�Ŧ�v?�uś��	A�p��V���Ҹ���%x�;��?0�����:������7Z�AbF�ߌ��6�a�{�t��8%���}75W�`��p���`�ݟ���o���yr�%ј7��6B�gjW�����ש�>�	2����lq\ީNvRrI��bb��=���v�0�~s��G�����Q5w��'A�d�I�j^
��/�	�/vx��!������e��jz�89��85��.L�*�a�E폄���0ixN�����Y�k���|d�h��JBbvӨ9rM$��[���^q^\)�|����s��9��a��T���
��\풜�w*H��ML^9)6La���h�-�Z)��&�� �'i�Fe����!�)8��Ǉ�-8��ǿ��Rl�������X�=e&r@Oy�G�����uz9�Ku���\
����A������	����H��+�1��Մ��G_vT��0�RQ)�˄��=6D7,�-wT���*�,z�5^� �J��.���������}\g��AV������������W���0u����0D�N�%�f�#"_z��|]�wߝ��hCܕ��_f-/�'dh�h�!�k��EY�F���/K��C�[)�U��g̐��9h�'�t���,�J+���~��X��]�������2ѻ�6WT�f��Rܥ��k" :E-T� ��O��4��z8�hG�\z�P���t��-O�xG�����>�ΰ�!��](`���{�i��x���9�s�_)��3���������*��ZÔ�d�4$��(�Г��sȐ���H��pBwN��[N�Q�m��~�j���<���C����	~;ӫ�\�粞��-svU}No?�덗���xE,(��R�G��戩S�@yލa_�(�6m��e|�B�1��C@��Y0����q^��c�������q��M��@��^�������"uV,$ȒR�MJ[3���T��J+�ᜆ�_����V�n�"�ϲ��K�l-���CR��X���:_�����]��^��\eKa��R�?Ī�Gg�1��q�p�\��@Qn��0�bNV���M�k����eN8�lu>��n����]�

-Y��t���Kt���P��q��G�M�5A��Z��xm� �>	v��2��G0ӥW8N,%5tRT��"�t&:Z�G�����V���r�� �U�)��47\��~~ү*:�g٘�L�m�:_17D�7D��$J�k<�V[3"�'L�J�j�c���
j��)c�oti/��Ph���#S���}�s���b�l0I�C�1��<FF��7=ǜV��O>�v����}{��#[�c'Gi���`� c�����|���a�
^�@��R:$��.����[��8[�T�*�@T�2�Sԣ3Y'--�Z� ���t��-X�.��O�5�E[��Y�1�,	�>f1�_[�ߤ�Єuk����TZ��1|���ɪMT;�'�҈�.�)�L�� �K-�m� aP1,�����������<:�p�_��k���sD��y�ѳ���V�N23�������̿ɷ�[)/�F_�,&>t2�����>T"�LW^q�������g�CX �j���Ƣ��bb�Ⱥ��I���qR�&�5O*�� CA��4�$<K��(J����轔ߴ���a��ξr<�ZvwX�#�ŬY'�y{�5B�3'9q藒��X� ��R�����C4����,F�8�=?�{f�hQ��i�>����,�a;��wQ4��_M���F��-W�y��W�7����;�T�\�=����c����R�b@�/K����a]oRj����[�-0����S݈X��[7
ȃ�kIy��h�O��Z>�?"9�=�*���e�f~���E��{S����[@@e p�����!��aQ�ԎҪz�ZZ#��sQU�^���Y}d��H�j7��M���R�i������QBp�:�5�_꼰Y��a�^�)t�L��{.xIN�I:�����e��%�[ԓ��K�r��CL���D��K���s_8,|Jc����ٗ� yB��Ĩ� ;x�	�@}�6Xw�<��%��	/����b7S���/�	�is#6��ǻ\Ia_SsF
ű�����X.�K���|#R�;�}S6�(,���/�v�cg;+
�����
E˼)q�7�E�h�}�[dبCa����'K�4�'�-	
����UM�����&�v��V�TŎ�iNh�{ A��(4�g4"aEN�|���*U������+|�iB1-*��w�@�c�16�cz�#�`2 �hì��|��ﳹ1���/�sy\���}6�u���Ygl�?�)1��bs ӭ^?6L���S8G��!�3�Z&�G:�n+���l�)�V�ī��`o��2��S�L�ot ��8�
;��]���3���-����Ο�T�g����5���Y��Rb$�sƎfQ6�a�P^����F�ըS���vӨ�S :eJ����	�V�l�^����<R��#��L�g��[0�v段���H�Ȗ�>g�\�"�_�����iF"�4�	��ק��Y��1M���|4�Ʃ��τ���{�-�+q�W����lX?'��}���7ި��Ź�AT��hHʙ�<�px�1B>Yⲽf��y��ԩz����]iR"nP�����/��@��1����ͣDυ/�z��7�L����Zx�S��Ҧ�6��+-�㷵� ��;���UZ����p�{��#��a�P��%�!���K ~C4�7��R�s٦7�Cu;�2�83/���A�Y�3R�����g�U瓙����yN��ܿFM���oF@��xu���y�ԑ]�Y��x�Jc,y��q3�����ƿW7��y���n')%o��v�t�߀��ϋꥲdZD�I! �V�2a�����8g���`tY<�'u�o�j�e��c�B#AR֏O�-ne0u�{��܊��g^yd�Cf`��ν��:F���+?�;�@�۷��_���H_�C0!����mg�Н�x��@��b�Z�r.j�Q8���^z|�߁p�ڷ���fk :��$r�`�������'vD�� 1�[�Kpr��\9Ҝi[�ErF��
9ҵ�%�~�v()�tc%H�ǀ��uB��_���T��K�� ��ؑۃA,v4stQ�Üz�3f<���F�c6�������!�2�W�+4t22�y=�o��u��8܇&W�ء��(��$9�/��@�7.{��u;���:�^l�L�5��P+p�
�IVe*I4))[�NP�D<���l	D�s�������1J?��S�)�Ϯ�jÖG��S�BU�)CtQ�����Gg�l�N�L���Ե
���7(�F�Fԓ��7�ƹ^^��٪��``| �ِ�n�鴛�tk�y����]��HzAf�\6�d`����/u��
�A
I�4�L��A'��͜4 ���v���X|��𬱱�1a��ұ7�3�e��|DՇ���´e�<�-Cǩ�b����I6�']�j�<�4�'K�B1�����F� �*m����w!��NZ��6�V�T񈍠��x��̃�9Ph�a�f�N�:l�ʋ�=Ћ=�2����V
�\5Ē_��<��Pu�J�@�*2q��okߪ�
}"���>mą���)��-�d���Us8 n��a\��x�.��s�?�=�
%^W���M�gd��r��huU��1h��4mI�M�k��!�i�����S����O�EDLGܰ���#$ u-h��0Y��wi��3���̽$Y���{Pt[Hr��a��S3��;p�Ƴ#(z �:��!H�nrߜ�$�rn�T���[�T�c5����}T=���o����������O���{��o��8~����2��k�t����z���c�^Ul�{$¾0sp�1F���,#|ݩ]��M���3.-Q�Р5.���������/u������1����7}]�x-�Pj�Y��J�G��w-�wG$�̅�
u��32��-��g��������ƀ�@����e�����Uf�;��3D��戾WV�id��l�廽~�c��b���4t��a�ә�d:rMֱ�[�D��M�B0)�ڴ��m�a�T�>r��'^Z}@Iٖ��s�ئy�ĺ"�Ӏ�����l�	cr�Kb^ƴ��eW�5�Z+�.�8������q곧s��Q�Is�#��^W�x?E���
V
�y";�)�~��!���q��	o�;52q�tW���I'Pn,ʸf���GW�N����g�6��8�����y��j����kJ�96�k4iެ'�p���FQΛ��se�Q�%��/�I$�B%{#l��v��A% ���U]�"a+I��&V��X�N�q��Nr����k�6��?��a[��BD�'�����k.���ov����\���x�a`����&M�m��_W���M8���`�ݠ�)%�������gSc��cwY��=����|g?�
_^
'����91q��77�Jx�M�$b4=Ĭ\>�?�Bz�����s�����T���U�mYD��J��+�΀� {+aw��jaV��f�����V�q��}
�0i�0�������Π���G \Cĭ�D��|��=~���}��_�D [M��X�p��,m�+���,QW>�(�)ۭ�`Y�	:W�t�뤁�`���VY���)o�-B �&�q[��%�<�>�k�C�I�_�=�C�y�V���c*�1f�XF}�����|c��4O����цL�r$qij��a�����f[�I�������z �7f\�H�|S�>+�K�_��*&]2㘑�m�?����������\�Ƿ�j� $�yּ�[����ֺ�n
m �������V�.ϟӱVl�T贰��Th.Z�µ�
`�4m �/$�Yg\2/��t�����ܮ�[AI��g	/���L��,u���
O	L҆ɾ��݊N�H}Jx���ᶞM�& �k�����+���kՃ���҂~�c�61�����0��97�2���{��ݦfTX����V�D'T
*cյe�C���DP�m��b��k��j�1.:Iώ�u��(<R W�ꡒj���x��?od0Z�Ƶ���mV�<`B+�5�dZ��<��mf=2.�n��`�^���?3�Pr7+G��|{����v��?�#˅�U×,n� G��z�N����k���qɊ��p������K�G�ʞ<�y�\?���x������P9�W�>��pk�}�~`F��m�%JH�B{�Wޝ�`j�����'��'u#2��1ڦ//in�&���x!�CrF��Z=�SN�O����8sχ."N�"a��:��ʶ�ޥɧ��و@��>eZ2��p�F�9Hi����ʣ���@P�>AC��u�s"EQ�`���z���D3F�C�v�3��C/�ϡ�G7��M�6�vO(����mY�x'�gA�ڈ"X�r5��)�af��B�a)�00�:����<A�T����,�l+����X���˸�'�ŀ��������F����Pf�)ii����+�Di���{�1ի��~�֠��Ե��9 �d������%)vJM<�� o/�ұB֑���T�ҵ�{1-��D��~\�U�^G�!i���Е~�e氐�8N���D��J]e��}�8f��Y{K��>�3P�z4WHfg$"�����D�!����%q�7N�LC�E&V�d��>�q�A8C����Ki��<��\�af�H�Y�u� �hq����CA�|���Z�<n�5Oz�>�%%$�Y5���_�E>�G"� |C��nw�{�]�i{K価���b��2��el�Doa&ԃ@qa���V�!47N�Rx�Q��Ks��� �����5A�u������s([�	���v�mΎ��@{M���{�g��pJ���[LR���W��Ra\MC6q����MxVe��\�^L�Vʄ\��o�.�e�5�M-FS�?�=/�4�TM\��u�\'S���z���oö�	�~Rsn�˗xhǞopk���_�S�\���M�Q�&��n,�$���8�7T��s
`�q���Ĥ��;-NsE'z���S�"��X>��q�͉�ɞTfA��FW�ͳm�.T���6�i�{V:�œ�.\�^��L �ʧ�F��[�q�/��%�L/
 �;�"�*@!�syL��
�����
����ܧ�`�=�����x��kJL6�7Ζ=��mV͆u�z�o�T�W0����hy�OFT�%G�^�c�̺~U'cw8j5�'_Y�n�>;�J��E(~,���Et���V$���\F�Ȧ�I�jl�ز����Y{�"Щ��C8S{���J��h暠M��ۿ\�����
u��/?l���@����B#,�;�>x������:b����$
8�� �16(�m�/��R	߽L���c��XBO{(��h�{�2"	V;��ou�4{�b�fZ���PU1&So�GlWo輎�*r�3+"V���i���3�K�fq|'n�Q�y9�w���T?Y������U�|97,�ޘ3A�s=�������7�w!��9�����FЦfI��C�T9TXI���%X�U��E�ô��֎�����~C�"�ex��G��vd�8'@��J_�p�I��ܜ���e�$�v�r��F����+���g5�t���qC>�pL������8[xiS��;�Z���f��~��u�c�� ��9s�%����MpA<�Z��g�I
�8>%�U`�t�p��(���~=��2�V��W���`ƃ�����99̡{r�@ѭy���.d;_�^{^±1��tD 뺔��o3}�%��I_�ty��C�?�|���kS:<
T��i�k�\�j�	����㔈�ӢG)*�-3'v�N]�A���O�Kkʏ8���<Z%qhƄ��r�`��Yrɪ�
'vw�찐��F���V�X��z؎؛�%�T��f�q{�p� SDX��Ǩ=��Ğ"A"}6�X�w��#��j�6
�����[$��������6�.�&hVV�Mb�?�O���Ļ�o��.�:�F_j��8�Q��נ	s�uRd�_���;���,��\��f������޸�����)�n!q1�,+i�}��ڬ�awY)�9�J�gv��着��@w�{���U�^�N��Ev0���*�a*	�EW�x9��\z��|Ɔ3� �x�^�2�0Pg�5���6v0����U�
׍
/$:���@�����n���Ca��A�MD�,=C4��}����qSR���	:W�XV3�- X7��q��b��ؔ�I�� ��d�Vb>a>���Գ�L�A�U̧>�Pْ��)�L;��
��궪Y��"�.�}L�,�_,��qv�<�M�]���2�С��9;���͏�x/������+�Y���΋�hțF�w�k;�)D:�����8�ܴ� �+�Df?�ez+�I+Y��*�>hh1!�D���{��[��5<Ya/��y{ʴ��k�#D�(c9��Kl�]�TGS����~}���>m��O�������n*+����2֖�(#n�G�Qt� qJ�gQ�B@�:�����9�,GD3�Q�a���,���X�}������wI�w.�AH��0��:5k�8���N�D6t�I���.�D<c��Z�.��Rd�9�jGM�=��I�<;�K����T�@ �oj���*k����QA�&y���W�t�0t�@o$�5��CP3��ts���f$��ۨ�zQ���D�Ι6���4	��hs�R֔�C��%�D)h~�HK�JN���{�,�	��w�hwy-r.S.��]s2������2"ÃY^}8͝YS=٤$	��A�Q���ݰˉ��Gn��ީշ�!rs|�Q�Tv����v�N(�.'M�Q_�����>,X�/�\K�K=�>8��O��c���ν�����$��GW\��5M��,쌗����J���0z��A�j�!2�m��?\��퀥ެ��B��u��^5�yb@K��w��ˑ���0�I4
qh�_E`6E?A�J�<�C��(��0a~�%��6O�@������kZ��)�&{аqް��1ZB���;)?�W��0�O��Oh.���bH�^����� `U���D7�Ũ�x��t�:����4�S�|V<LM3����_��Xx"�I����{�DDv��]�HV��^�(X_�1�3-8Ϫ���x�����~O2����n������/DJ�&i���*��X�f�r�i�����=x�-&���ҝB���d��iD[�:�����BF'����t�ߍ��ZF��qGh7ؓ�/N#��OZF��Ng���=��SL��=R�
1�k�@W	C��^�&ׂ��-�����������*2T�zN� E���N����8F���B��� �>��
�gVh]L�u��^?C	̶\Z�'f��p�C��Z��c/I���Q��CC
$���>`�w/��Ԑbm�hs�7R ?�6���ٝk�ǥ�