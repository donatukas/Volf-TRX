��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~�f�?|��Ť6
Y���#�J�-�k-@�*DE����tF��鐷o�s�s��o��kۣV���s������I��`�V��M`�5�~M�8˄7{v �������d4����S]V���0lm���U�Z؟�#c�.�X�ȡY�D�~��K��2x3�mlk�\k��zQ� �����i�4����k\ k�Mg��y���٢�N|����� �U߭"��AZ�f��gDL0���mV0�y����;F�����( A�:�f��⋫�Zt5�(mm+��N8�.uϪp�-�kAt�2�?��Mc�t>�nȓ�{�:�$���vB
ߩ*.e�Ɗ6�Cd篓%�+��М�Oj�Ǧ��x�AǌE���Ki��v�X���hk�M��P��σ�ﻖ��=�Ƣ�Aj�N��'�>-��GY�H1.D����|�%ϐ���ڽdTV��nU"/5���Ʃ�;o�h]W�8 �<��VD�:��Ɖ���Yc�� Jp)@�,��8�%<�����A�y�,�Q�~ [�x��M�C�o;�I�hj�t�J�1̱���ӅG->C��x%�%�+&��b�N��e��x�Z��^���T��Ef��^�c։W�7�����
��?��to2����ll�ɓK�%sV�J^��0~D ��ܒyBk�I'�4ߌ�l�xv�&;�u�E���'i��@nžm25~$���q�%{)O*�*E�����e�MsF�u�$��_^|��Q���1N4ذ�b0��!Z,ӕ�^1*G	�fR��~
Ie��Q_#l��Tgr�K̾3��8CGRd�Jrz@�J��&U��a�w��9M.:���0z�!��,������V�E>��+�-�w!5%�n'�j�r�M�%2t"���Ŧ0ĎY���~��TSX�����Q7��\r-��x k<{�C�M:����k�m�kX}7?e��-v(n�������k��K�[c�z�c�ZD��7N����ף�O]�W#����Fo[J�&��.�[]�uE���s�פ��+>#���]�Q�k��2�	�@L#�7M�*���w�i���#j~ K�2�rl欢ψu0,Dj������]e�=nK���2�j��V&�J:���e&
qj������gN�ec),(��#��_�a`c������Y��篶<
4���m�+N���m��˝{jA��r'���`�`�Y��p%Ly�'���Y[������LW����=dc�j-�s=;�|�k|ѿ6!|9������D$[�S�ɉ9N��Q�>+l�{B QP�%�!����:KW��;M����Z�HM:>��}�t�äS{�S!��J���&'>̤�%������y�k��A�4�bz��UH������4�&��|�.tQ2]��OR�S��O.�1r���V���jĀh���a���k�+�^h�V& �Sq��y���-bj����BTc*����_c�J�I��V���3��=�BdY�쉁M���) ��\�P�g�*0��Q���脄]{S�$�qj�l�֛��xR/l�\L�$�v��7��~D�`�����gG�����c�;9���b���y>�]45W�X�������X��5N��U�,�xx����B?��b��d,E1�|�įf�8�p	��&%���4����ɉց���_��f��u����Z�N	�xeZ�:C�:��O���X�CN���)`;Ol��Ѕ�P+�bOp�/I@���3e���������!2��Yx��G���\\�T�ߟ0��?�Oz�|"z8U���Q&�Iw{�4W��HBCȎ�N�Zq��"4��|G�j��c򎟑b�P���]&�EV��&E��5���R�#���ۅ~& ?���z'�0�>��aW]�h�8��'�LF������>t0/�(�Y@
Q�+�����)�/���Q���>�]|��afY�����4 j���d%��5ka<��XС���1�F�=�7�o�$R�u����
� e�� ��Ϸ1�����⧇�l�?#����
� ����S�G
DD���e���K3
�<����tg�ǲ�t�k�X��+"���<hՋ�秼d���3������.��u�>e�	X�~s9��;=J?��dl�ρ�P@��=>�lYs�L�2V�,�A/�}���c-h�P��pS͹�ך�ƪ)���A��\d�W�Ƒ�j����.�Y4f�v�h�'.7��_��9�6\/�9��([N����������-E��)n��FIX(�� B�\z��! 9�G��{Hi@7o;^�	B�# �^��Qyf{t8+���Jm �����)Ӆ�>��w��gP%Z2d�v�(r�s�NF�a�/O���ګ��KT��O� D��ԟt��&�y���8�RgZ�!SL�im9��J�F "8���-�q�WĀ|���̣w,��D�w�=�;i�"fN�qk�)�%�Xl�,����y�C��i��sK'��'�&�r5� �s_.ġ�����T��ϥ��qx"/��mKW���ي�k�>��LסP}����P
�MF�Y�\)O�W���V���:7�]_4t<[�,�|�����47/�62#go�c*Z��o��L�I]�E�ʼ��|7�RS��Ʋ��	�%�)#J(�v�Fҷ����|��Ҽ?)S;�h:��#��N��c�+���>N
Ԃ%��3˗Q�������zk;�qa�ׯ��)f�&z�kɊ��trT�DX�ky�,}�o-�e)��F�Ilx5B�֐/�Մ��Y^���U��P�����Ɨ�x;��u݅<��x����