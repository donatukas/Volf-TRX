// megafunction wizard: %FIR II v22.1%
// GENERATION: XML
// rx_ciccomp.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module rx_ciccomp (
		input  wire        clk,                //                     clk.clk
		input  wire        reset_n,            //                     rst.reset_n
		input  wire [31:0] ast_sink_data,      //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,     //                        .valid
		input  wire [1:0]  ast_sink_error,     //                        .error
		input  wire        ast_sink_sop,       //                        .startofpacket
		input  wire        ast_sink_eop,       //                        .endofpacket
		output wire        ast_sink_ready,     //                        .ready
		output wire [61:0] ast_source_data,    // avalon_streaming_source.data
		output wire        ast_source_valid,   //                        .valid
		output wire [1:0]  ast_source_error,   //                        .error
		input  wire        ast_source_ready,   //                        .ready
		output wire        ast_source_sop,     //                        .startofpacket
		output wire        ast_source_eop,     //                        .endofpacket
		output wire [0:0]  ast_source_channel  //                        .channel
	);

	rx_ciccomp_0002 rx_ciccomp_inst (
		.clk                (clk),                //                     clk.clk
		.reset_n            (reset_n),            //                     rst.reset_n
		.ast_sink_data      (ast_sink_data),      //   avalon_streaming_sink.data
		.ast_sink_valid     (ast_sink_valid),     //                        .valid
		.ast_sink_error     (ast_sink_error),     //                        .error
		.ast_sink_sop       (ast_sink_sop),       //                        .startofpacket
		.ast_sink_eop       (ast_sink_eop),       //                        .endofpacket
		.ast_sink_ready     (ast_sink_ready),     //                        .ready
		.ast_source_data    (ast_source_data),    // avalon_streaming_source.data
		.ast_source_valid   (ast_source_valid),   //                        .valid
		.ast_source_error   (ast_source_error),   //                        .error
		.ast_source_ready   (ast_source_ready),   //                        .ready
		.ast_source_sop     (ast_source_sop),     //                        .startofpacket
		.ast_source_eop     (ast_source_eop),     //                        .endofpacket
		.ast_source_channel (ast_source_channel)  //                        .channel
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2023 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="22.1" >
// Retrieval info: 	<generic name="filterType" value="decim" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="2" />
// Retrieval info: 	<generic name="symmetryMode" value="sym" />
// Retrieval info: 	<generic name="L_bandsFilter" value="1" />
// Retrieval info: 	<generic name="inputChannelNum" value="2" />
// Retrieval info: 	<generic name="clockRate" value="61.440" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="inputRate" value="0.768" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="read" />
// Retrieval info: 	<generic name="backPressure" value="true" />
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone IV E" />
// Retrieval info: 	<generic name="speedGrade" value="slow" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="-1" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="-1" />
// Retrieval info: 	<generic name="mRAMThreshold" value="-1" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="reconfigurable" value="false" />
// Retrieval info: 	<generic name="num_modes" value="2" />
// Retrieval info: 	<generic name="reconfigurable_list" value="0" />
// Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
// Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
// Retrieval info: 	<generic name="inputType" value="int" />
// Retrieval info: 	<generic name="inputBitWidth" value="32" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="25.88184,-11.77676,-42.47139,14.62374,64.98443,-16.19333,-95.30045,15.43182,135.7651,-10.75484,-189.2556,-0.1792373,259.1529,20.65105,-349.3771,-55.22246,464.2181,109.9167,-608.3312,-192.6859,786.347,313.5165,-1002.837,-485.0395,1261.6,722.4344,-1565.65,-1044.216,1916.052,1471.749,-2312.049,-2030.281,2749.287,2747.798,-3220.302,-3656.454,3711.905,4790.396,-4206.394,-6187.838,4677.782,7887.381,-5094.268,-9931.155,5412.869,12358.98,-5583.896,-15213.26,5543.345,18530.1,-5220.412,-22346.94,4526.717,26689.58,-3368.222,-31583.84,1629.933,37036.99,805.929,-43055.5,-4081.676,49618.68,8337.356,-56705.22,-13741.61,64256.33,20453.14,-72214.42,-28664.35,80472.06,38547.0,-88927.47,-50313.76,97413.95,64142.51,-105778.5,-80262.79,113784.3,98851.55,-121220.9,-120154.0,127769.4,144340.8,-133155.0,-171676.8,136961.5,202326.3,-138839.8,-236587.8,138251.3,274629.2,-134753.3,-316815.5,127640.2,363347.4,-116332.9,-414724.2,99869.66,471247.0,-77438.17,-533684.2,47634.23,602587.0,-9184.515,-679272.8,-40179.41,764883.5,102762.4,-861920.0,-182757.3,972972.4,285110.0,-1103365.0,-419068.4,1259662.0,597716.7,-1455176.0,-847254.9,1709824.0,1214643.0,-2066687.0,-1812364.0,2608282.0,2938129.0,-3544861.0,-5781064.0,5218750.0,1.94578E7,1.94578E7,5218750.0,-5781064.0,-3544861.0,2938129.0,2608282.0,-1812364.0,-2066687.0,1214643.0,1709824.0,-847254.9,-1455176.0,597716.7,1259662.0,-419068.4,-1103365.0,285110.0,972972.4,-182757.3,-861920.0,102762.4,764883.5,-40179.41,-679272.8,-9184.515,602587.0,47634.23,-533684.2,-77438.17,471247.0,99869.66,-414724.2,-116332.9,363347.4,127640.2,-316815.5,-134753.3,274629.2,138251.3,-236587.8,-138839.8,202326.3,136961.5,-171676.8,-133155.0,144340.8,127769.4,-120154.0,-121220.9,98851.55,113784.3,-80262.79,-105778.5,64142.51,97413.95,-50313.76,-88927.47,38547.0,80472.06,-28664.35,-72214.42,20453.14,64256.33,-13741.61,-56705.22,8337.356,49618.68,-4081.676,-43055.5,805.929,37036.99,1629.933,-31583.84,-3368.222,26689.58,4526.717,-22346.94,-5220.412,18530.1,5543.345,-15213.26,-5583.896,12358.98,5412.869,-9931.155,-5094.268,7887.381,4677.782,-6187.838,-4206.394,4790.396,3711.905,-3656.454,-3220.302,2747.798,2749.287,-2030.281,-2312.049,1471.749,1916.052,-1044.216,-1565.65,722.4344,1261.6,-485.0395,-1002.837,313.5165,786.347,-192.6859,-608.3312,109.9167,464.2181,-55.22246,-349.3771,20.65105,259.1529,-0.1792373,-189.2556,-10.75484,135.7651,15.43182,-95.30045,-16.19333,64.98443,14.62374,-42.47139,-11.77676,25.88184" />
// Retrieval info: 	<generic name="coeffSetRealValueImag" value="0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, -0.0530093, -0.04498, 0.0, 0.0749693, 0.159034, 0.224907, 0.249809, 0.224907, 0.159034, 0.0749693, 0.0, -0.04498, -0.0530093, -0.0321283, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0" />
// Retrieval info: 	<generic name="coeffScaling" value="auto" />
// Retrieval info: 	<generic name="coeffType" value="int" />
// Retrieval info: 	<generic name="coeffBitWidth" value="22" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="31" />
// Retrieval info: 	<generic name="coeffComplex" value="false" />
// Retrieval info: 	<generic name="karatsuba" value="false" />
// Retrieval info: 	<generic name="outType" value="int" />
// Retrieval info: 	<generic name="outMSBRound" value="trunc" />
// Retrieval info: 	<generic name="outMsbBitRem" value="0" />
// Retrieval info: 	<generic name="outLSBRound" value="round" />
// Retrieval info: 	<generic name="outLsbBitRem" value="0" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : rx_ciccomp.vo
// RELATED_FILES: rx_ciccomp.v, dspba_library_package.vhd, dspba_library.vhd, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, altera_avalon_sc_fifo.v, rx_ciccomp_0002_rtl_core.vhd, rx_ciccomp_0002_ast.vhd, rx_ciccomp_0002.vhd
