��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����E�"E���[��D��֫�>���B����5b�$GK����r�
A?'����%*%���C��Y��g
�3{���I�=���M��fXr=��6���2[��/�u5K�<��歍�ιk.4��0i�]�
y��]z'��XAh����˟�@�P����_SHIC�8v��9�*�iv���[C˛�:0hR��N���sΨb8H�kt��EOw� ��i�8��m#��<aF8�����[��p]2�=3�УQ�k%���>k��
^o&)��"��D�5��$��(���9��h�&��|�T!^:)���'-��ўg'�mD\i(�vn�EPM��|��X���jխ����vj�إ�mA�����ܫ�}��U���YJ�¹�{o���5�-�<��N�;�k��3��PP��`���n�3�q�P�ǜ���/���jx̛�/�Fq�]Q���I�J��S�N��y����X���#����$(kDF�~Ʀ��P�F�l6����á�v:s�\�P�����1�<�l�x���l�xvo��+;pȎZڒ�[����I����+�����TT�-���mb�]@�������@3���W��5�F��|�E@��5���|��b�+�����ө�=��QW�!v�Xw���KQ(��1�w<�n�F�Y<�Z�҄6y��!�y0am�����?̒B�	�wO�g�#m�*�3BtbT�[�܉` Ƥ/Ȃ�b�K�v�^��p�+^��p_�rr�'C&JU�K��1�jR�S,������v��Xh ��u@掶v������r�6>_`��B��2eG�&RUC�<nROR�OTqa�|�F'�Ɖ^4B1�_����g�5�����5�y��7��S���J�M�����t������j�9�U>�1K��d7��Ώ�0Λ���8͢��7PS�@���`x��9Ts�Q���u��^�-x������Ud���ۓ�G�#$+��}�4� �����6��9�����`�_����5���Z���M�0��C�,W[�s;a�b�u4���5�'p���_ׯ�9��s��ޑ�j�W��_�m��V8�||�r^�;W�i0��I3x��	3=۵�� 3$�c��/�h�l��AW�:,%)�A���]��w���0�r;i[p+�pr�k�
E��$Qa8�m�H�H�*�Pe�8���ڃ���Y���4z�Y܏L�l��P��dx`.�J�F��|�&�1y�������D��q��s����%�y'� ��z��컎�v�f�\�終`�]X�-���S�U�536��%�ҧ�w�1[�n��X����j�ض͑s@�����l�b�I�_)�o�K73��td,���I�� �+ �a��� �RZ��[@�X�፠���d��ј�{ˍ���Ԇי���8<�C����4�:�U���b׌�cn%�o�q�i�$��9 ��ͷ}��j��� +���X[]�U�R2i��ӧh���"D"���@>.QP�ځ�	�Գ;��j�M̰�_��Y ᕼF(F�ۖ�ss�<�J�&
��E��_��ێ�IXO��@?P)�eMa;�|��w�[����Ԙ���G�yNfr��B��@�89�
��Y�5`�4��+���:8M��|�j4q��WӦ���Df����#ȕ^������(Y��1��I)E���� :sJ@��D�q����b��W��ϑ����\ܷ�˫��~�g��3ѱE��E��'p��&`��fH��*�;�u��C9Ҿ<w�q;�k|���(� �7��1��9�y_��bN��Aː�@<m�S(<�����z?��m��zݥk�ʐKNSN�<*���"�聲�q2l�8�mL�K�r8����09\�zP^����I���4��Ͼ�tűr��jU�'+C�c
��+%zy�D-��f�Q� ��V(�4��ہ�S�(U�D�3�l��5TRH�Ǥ��7�+���K��(��)K���l��ZMg Nԋ0 �r�zR@'Iϐ��P�y��\e'^�)h�!s_�]� #f������������4���j?�y��&Iܢ�p����K>J~��Jk����j�0ܩ�##};e_vB�8_�jD�2�X�2W"zONiS�%�1��;�AX�!K�Rv�$C]@��cŶ �z��4Fd;��d[ L�%��`r4�Q � u�F�p�՗�b$��3�:A)c�J~�j0��g>�eG��=l�����]�4�'�ߝ����c�-V�H��nc�w��^$�����ܤ	���"��^�T�>�z �t�:��awa�GW�6(�?�2��Б��93�8D��N�y��v�d�� ������u�⛻�K� ���&a2 j�u37����%�X�ɠ ���O� G0���q��ӡ�w��o�h��?$p&|�1�u���D�cI�;�H1O$�ϴ�>��=K��?ƕ�Dc�Ȗap!��?�3Ol�����o���m�Ŀ���Aq��>��*6����L�c�m�EJ��'hKy+xvGvSD���R��}��h���#�*yW�+�;�����R���}xe{0�5�7�w���� �V�=���ByӃL����t_W]�Q��q����b��J���* ��5��8�L!D~X	�&UCѧF�p_��Û�>��&�X�|�]ճ�Krb)w�aت��	�<�JM
)�	?B��OsA�W-�RY�3���K��`�>5K��x����X�8Ex2�5����J!��#��׫͑����	��*�uծ(��enJ\a�^f7iƝD��	"�Nu�a��mvR2i9ď=�皫����U�@@�9�
�'����0S������*!,��/ui������+��H�V�ePC�e9��n�y:,�)
���c���;ӌ�Gg��6��5��<���p�����s��
68�`��E��k��=&�u�S��p˴��~�s� �!���\�~�b"E�D��$�"�z�K�v\��Q!�d|�d��Vs�0�]��jF��{w���l|fM8}�ra�PeOaS5���	0=�J�a���OH���M���E����x���8�8��l���+]%���]�Kt|�A �iu:�o���3c��lr-9ݥU/![Dd�E#|���#� �D�UX�o����hn��ӊj3P�8�~�,N�C��k+��	|�Ȥ�������F�0d�\�W+V����8E>s�1�֧w������/�}ݽ�Ȑ��-N,o(��0�{�A���3]+��P�HP��
����Y��U��Ui�v�d�^D\�x�s��о��HnE{#+�,���)1��{�'�l �.
ﲑ����+��?!zd�}�uo��[�H�����$z;@�Xg�A��1�z���NV�(��U���p��,R���q}'���v�8S6'����U�Fb�}Q8���x_�Y�-vq�"��^�7K\R�&�5?}eZ->�?zD���tS�5���N��^\��@8��s��֝Wv檃	�鄗+-p~���,]5���k���ξ�F��a{�xƏ�O��Q��A\�$>޵Vzk�ڰ<�\d����3ًk�:ǧ���I���x�m�!�����Z)���@7%�u>T���d���Ղɾԉ��&��^�l?���j`hH�[tw�N����y׍+rL��iu�r�����X���84$���G�����-��C��@�m�ګ��N6S"R�j)�FQ�Hc���D|rX��͜�e=��u��5ᔻ	�j�fm��yЇA{n����R K�����/�\�P�K�]9�\Ymr!h��r��i�� �\A��S+�dR�,>k��J^��'�bT��]V��B��}��Խ�k�D�I\�v��g��l}��s:��7޷k����0͖����ɛ�o�* I�R�hQn�/����j����d�m0��8a~��,r�����Q� �U�1��㤸�F�;�&���:��hJ)[y4�M����I�=�u'q�w?4�j-&��t�X�$54(}y��gs-O}��_�� �7?��J6z���i�'sHo��LvqGL0�z|b{�wl��_�'3�Z�r(��o�δŒ��>"ћS�F�)�N��m��}E��?4̰7plT��H9�&K����T-���vG�����	��!-$X	�T� �OC�=� u?���j5�}x_4�]��Ko0�"^an�FS�z����/?�5㢣�mP	<S�B�Ֆq��9��yz�6o�}z��cx���HN;C�����a�U����'��<;��(�U[S�d:V���=�+��OhB��J�q:`�Q~/^fF�3o�L�"@^�R�'<%||