��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.8�KoꃦW�Y7�RڦX^���w4�N�E�|�y��xJ"F%X��[DL��TKg�������������eKj]���C�����̌��%��{u�~2^��� �L�-�)&Et��Wu4��ΩЄYQ�qh�.[̽'�@Ɉ��v�H�`�J����͚)����י煄�X�z
�x���W�����4���@���Tu���^�ҡ6��8!�f~U7��jv
υ�J��T���
���f��(s�r�����"���2��ǖ �;�j�^@%үD�����wV��P[�q;�C��N�t�9ˁr�����w�ܕE ��_}ZA�;�Y��C�p	w;�#��~�?��Nt�`�)m�|LY�I2aw�ϊ(g_JU��9q�2(Q���C�;hyJ�q�j,�]L9`�,�u�Q3�5<P��DQ���D�	��V�N�訛��|u�ǢL<\���X�e.VQ�H/�-���~��hMW!F,f����"E��A��Fo������"�Q�2�jI���^p���T� �!�}4��1�DF�U�� T�`2.7}��>��f�7��v�1��~A���6EJ�h8�(f��mjC�y��۴'��k䯌��}ⴋ��׬�W���ˇǇ���T���1(��/#h�ɦz�0�S��o�Υڰ�;�l�2�mQ7X�0��Oc�s\%7�h���(�K$P�����S
���1zu�U
ֽ�nY�Un��,�7���,��' )h���1���qBV�{�|L�@T �|��[go�{�1]	��}RR��)2�\|��~����`9<4�q�(�r8�0f�fx`�5 ���@x1C�N2tEO�fV���&�&^}�+#+�j�٪�Dݾ���f����Ǆ�4*N�	a)Z��\�V�Bi+�X�=��U�uZhk�)V80����!�j�v������=DJb���� %hh]{�if����y���4���Cso�;I (��,�<fYfˮ;Ecy��=d>���p����;v�)X{X/c�EnͿ�̙�O+��md�	_�y�ZJ�'/A�Zv����~|��8�K{g��K4ߕˋ/��D�϶� W_�M��_�%{n��9��}��w�;����HEp����c���'b�x