��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.yu�=�6Љ�u�J��u ʸN!�݃�!i���=�F{��މ��zM�Qܲ�gu�"�ӵ�����Hju4HG��PY31�����X�p�u��S=_��k�&�����*��Ӷ�P�,�S���)�q�m��B
&b'�:%T(e=Z#H����GV�A�1	����g��.r� �5t1�"��,�?�!����Q�K&ӣsF�O�S*�A�<�Ԯ�h>�@8���; �[��-���e&$�t}7 ړ�*e������H���rg���_�s*Z�K9��߃��"�]�|B�V2d���?���M���&x%��qޓ�Y��J=_�έJec�u�s5q"� ��鶬FCq=G#�X "$4vT����d�����̪'p#k�K�TS��0�CW�!���p��_*f��9�MZ,/G���۞��⅖%
.X/i�x�55aΎ}�.��݋'�
�ڴ�<`W�&��/9���V�G�l0���K$-*�_���d$��{Rq\3"�׼��s�?q�y'M����遼G����.��HkQXtx�+�r����*����ڦP�Ƞցrb�3�c�*�u#�j�g�5���f���C��b��6�O1��i(>�3E�w��J'$,/o�X��ʲŴV,_��<sz=�{�|�$xy��}�6*
�ZܪW�C�7�)�j�#)�$H��?'��7"[K2f���/��X��fޣ�r�E�K�;Cs��\ܒ�կ�)�Gϒ���DQ���息��6���9h�r���3�s	�C�Y��Jrz��v�=�p���Wߥ�g;(4t��Q�W��0�2�"W���V��sSL�HU�^�izg��f�0�֍�O��
5�����i9�M��Oȧ���ֻ;���D�^�e�dw_�pl���$&,E�ʕ�ާ��c�M��������@I������FE[ �ɗL.��]�.��_�=��{�6�XwXe��$ؽx�������������j��ޖ�|н�( Ȉ��I@\SYՎ�X=�U+��F|R��r��v6GtZ�7��I����2�+P��%����b���L�'
$9<|��PY��z`O����XE�߶��V���x)]v�.���>��B!=���خ+���]D�-����"�I�-�v�N_�j�W;�s����S�HlmD��&��my�7�����y��<Ӑ�J��">AS�; ��ft���(��9��PN�#�&�H;m���&5�i����:�L|S#�D�M� Uu�ﺔ~�5L@.�X��5����,,Ꜻ��aSIpv�9\_�d�mצ1߇�g@b�]ӭ�]�!^����%6q�	Aۢ��B"��<M��]^���Q�>�az'ڭL~q/�}zgQiy�{�]����n�w!���aJ�N��8��n�N���(�튫�0��#xT���f@n��񾀐)~Β�>�76	�m�G�R� � ���\e����bH��p�GV��d��NW��g�䅂����b�L��Op���^���e���&� �O8v��#'�[Z�y��/���b��A/�SD�/���s�g�-N���m��M�.�|G.�a�'�ɽ���z֜�1iE�2)Z��_%�:V�y����� 7�����YK)�M'f�mb\#A���-����T=�zG�ZL�艟;��[����0��oS��|NZ�Li���R�ښ�����Ge���𬦕�v)0��*�s)��+�pC��uN���L�f������k��8�t�V�>l�ӑʗm
3 Jy�_������K� u����Q[��M�J�|�A�}XV�{������C@�i�y�����HǶ	��:��8��m�ޢԾ]MۺV�7bZ�؃9�Z4@ɊXe|�^FvN�;�x��|����j��C � ������˙b�U�hE� ϑE�鄧�@)�zNا�Ti] mq�O�7�l+	���t��B�FMe~��ҫBgk>d���0��6ɣk/ ���߹�A�qs��ae銜8^	=P�]��]\f��JHt��V�H̉!�X�<	a�|��Mk��̉i1e/J<�H���.v�q�o�
L,qy�.��Z[4p���Z��1���h�7��K][�L����Ԉa���^�y�n��΅��a�T�i� P�Ig`p��@u?8G7W��%'?`�z�ćs+���΍�
I�L�%B���g���
�%��w/�gj�JOw�%Rү�);H4���zZ���UHG������f;_)P��B>I�f�����o�D=d�W��頕�	�OX�4m7�	�<̱�i�����4�гr4
��.�$��Η҉��[�х���J}_I2�@�7-��K�^p\�
�=��%�?o��qɰ�gaC��0���@�w�,��%~�*H}s�~�K`� D(k�d~�S!wW������jU�L�,1��el����6]j5�^���T��]2�]��G�L���Υ��A�ь'XkcЃ�ݶ����6\?�D���ڿ�^������bX����w)9_,Q��m�L�I�i�f5��D��'�P@V�Űgi�H�N�����}����/�,��V_�#��9�e��?Y�"�����icq>�ubbS���\�f(�l�_��T
�\�
�a���\0����~��i�#��/�*�B�y[�?��n�p~���`E��b	��̃�>n�n�+,B�C.m1j��\�'7W)6�ۃ�\��%c\Û�o5�m�t�i��G��)�T�������e��Ln@��'^�Ǯ��D����'U5+�{�E_)EFj���o��H�ʵc��A`.
C=���]��^�
lO�-b
�����������%�v[��]��2\��W���y�Ş��2��~�1�ݖ��C_ 4yݙ?##r33�_�#���T���B�d�[qeVp�Y�q�6�d[�,�&�'��f���)�Ga��&x��5{�,ǎ%#
A����nA�oZ%y�@/��s�8���3?+Mu���Q�����ʉ0�Vv$���Ն����BMnF��?�ד�cB��D�=a�ؾL�bZ����B��2Rñ���h_�F4�t�Ne���蜨��r\�0uD�1��A�sr欰�����vH�6&��a�Ȥ�xǲml�WN&��bA�ej�*��x������Pm<׏���}'.4��F؞���3�IT���n,�����E�S\B�YDs�V�$�h�`�������ɋ��H_���Q�5Rx�y�k�L����1�	����6�A6!٪��������Ֆ�*��[� z�%��αO��U��S)��ﶤG���i��;���<)�wr'	�e�b=���2�I���<�*� C�t�"Hu����Ĳ����^Mt�β�c{�������n_a�Q�6�B�8p��;�[�{�Q5;�;��(�.F[Y�σ��\J@{Ε�-$ۡZ|Swev,f���޹�t*Xs&��j�,j�
�����$�6mD�Z!�����㯀G�s�콼{�c_�E�	ǲ��j���:�r~�\�'"���eU)`��T7D�f�g?�bJb�H�"e5zN@�8��A�jE~�&��L�/We���G�(^��U���
����LJ׿=�#��U����|��p�S�qV�6r5��'��BF���B"yO�cGAF�4��yisȧ�
��n���T��޸��+�{�deVd}�~~�)���`��:��'�{ʿ5l���hf�I �i,�ə�K�Gﰀ�[]��������M5����X0��]4��z�Fo����D8�,0ԛ����2H�����~p��ɧ�������b9Q!�*w����Nϧ^��T������V�z��v��=�)-�#�ُN/���`�n��k�{�p ��O�����_L�>�	�^�s<F�T�5mOt����*M�`�E��7�0-
�(��U������8��W�nO4����%q��/�\8(���U��+�/�k��K�� ��Gwu 	����*7�.��r8 �{ezah�5KQP�-�!�ǚG�h�s�����d�åe3���c�^H�u�M ����Je�%�J�������R-8=�3*� �v�7[�������4OW���2����si2ព���B\��Zj�~���VqYf�=��ͽ�;1�h|�'��N"�n���i��
���b17g����@��~w(
�X�o�����q�r~-�m�Z��v�䈄��EK��$��-�p��l���ޮPq[]~�׃���d�����hj�r����yB����\8��H�����Uh��BE�:0X�Y{��23Kb|��x�P8�0|X!�E�`(��v:e��~yg��ٜO�9h��ӪG�@��Z�e�/�ǟ�g�顋�{�o{B�o1�ZS��cy��bNu�>=4H��,�76�l�Ol:�7�T���	��V"1B}9�#5�Hį�\F:OPA�qT������)�ܰx������ċ���P�?�pO�V#ln��F�����F9֛U❊����T��u��_R�jc���Cf�[��:F��Bm��$Rw�hG%�����l�=��V��Ţ8��x�G%t_�`K�sx�`���mw(z�R,(�Vn
�&�p���e�<jm�F�Cq^B�MF|���?���óGV�B�� �p�u��"O"�]u�_-`�Y!�=P�H�����6���Bn�(�o��U/�)32�U�M���oIc'�;�i���5��4��c��V��R#'�� x����aq�
��g>� ����k�X���7�2F	���.���(ѡ-
JM��30S{1�������A	K*�I��b��R��y	*��l���Z�p �?#g9>�=r ׉����\N5��A���E�FF���/me�!nШ���|�)8�F�:;z1�DR\��R���_lvx��8ՓB�dܐ�?=ɟb��P��Zx�a*��~ųJ)˱�^bWMc�}�\o�.u\�(fW�#��4;�+Eʉ1GT�4Ob�-���6���㢢��R|�̤���������ɝ�/FT=����S����� ��Z~=�$i������D�,�8B-(m��4�t�vs� �) Yj�Ԏ`��n%�_��#'��d�%����|���@�(>��^���b�5Y�_ß�Ϩ��Z���s���A���O!Ƞ�ժ��pZ����em�~��<��%�� �d�>��G��޽7{�m�>'�P �"�ŏ�V�Q�Ֆ�gh��ج!�Je����� �-C�EX�ɦNf�sԛ�(��J�"�rA���l��\�z6��.�=��7ؗ�vj�t��a�/��J�p��\���*P¸Z)o/SG]�.�O[��tZ�\�`�>��y��*���FIOx8���/#3~(��Y�����I5�^�c^�WJ��D,;,��U�������&�V��4%E�"�>�C��@K}��w�Q�6����%���b��6��]�S�I�XW�@���
 �X���ws_��*b�� {�ze͓�U��D=����U'(ߥ;�杏��-�t&�h�Q6l�^�NO�!C_��3��I������3<�ꤦY����K�'`�Ќ��w.�.���YH��@�[�=o�����&�}n�s�H������K��R�
R�x�!�u��;���y�	JX�(��:�a���%&e,v-L�7�/�Q<� D�8�߯#s$\'x�T�w�dcC�v�8��oR����Ě�&D��q�y���� ��S6�9�[��ށ2�q;\E��t�9L��qIE����0��&��8y�)]x�UbO����Lh�NR��R�o+��\=�)iE��o��v��<�-Bt���;m�m
$a�P���a���s��{4�U�*W�)���T&U����1&F%#
�[��1�e �ܛ�.!����BW���>=��E�vԵ�r(�-K�u�p_�2���c�B�֩Ͷ�D�]�7�3�	S��$}v�z�~����~��*�Oq��Oȟ��YI�1	'�gP��e�(�3�THt@�H" ��@S[��_*}F�=9!R���$5�U$%���s/�����O7݈�v;'�6�Y]%����ű� ��ky�D9p��R�����n�~����e��ey��Xh#(+C��f�Um�#p�'zj� W;���A*I�M���ɚ}�Vi{g'�έ�X+�C���V��+��#�O��B�G�Y�f�_ h��9g��U��&W�P^.ǧ������1aO���\q��U�*;]�A�{�M���>��\�m�)���R�y��,�nZip���G�Aix����Zi-�[�-��|�0�ܱ#���&P +���o2���m�B�>�f�vl�������<VR@�V��j�0.m��D��m�93�0l�׆+$��zI��{,s{����%���L�4�Y3v䦗��A">�m@�2�d��-�}�C�3��f���m�!��|H�RMX�b�:ӾoɜL�mJ��+J5��}S�õ�ޒ�PƳ�fk��纉�t����\�ׯl�U�����0��?QZљ��7��-ς�uV��)���+TPs�y_��yG#���Qz�>M,jr���;먷�0��q*8V "V /��Kk<�ޕ�Q��p���D���w�bK��Q�d�K>ډ)4�|���m�~Z]0�33+�)T�+�[���
���g!�[7�@�>�%���U�N������AHgdx� ��8M�D7F9�u-���Q 3(p�o _���L�\)�G�VB�T[Q�����c�]+"��ˆ,�wX�}\�]@��G�b	�<TO����vTlM��^U�=��z@�M͖1;�AH9N_ۭ�5�o�5�o�H1������p�3��d�.�.W\����ܱM;� �R�vuZP�!�֌8#���Fn��)� �3Ů6��,�s
M:��8J�=G�f�kmk�3|�u�5��K��壠�=T�[�I�sd硕��ݿu�a��,����&Au����sFq4��Xlj�mnژ��C�կ�I�8u29�ώY� �FF��E���+,�>��vץ;�i�S��^ �/�)I�b2*�b ��	�g?��O��I�=r#�"!.�����t&J��ﲣq�>��W�W�P�1���� ���KG<�R	���/J�dc�a%�[q���>�]I���jһT�i�j���z<�t�K�ѳ}�7e�\;R�V�;N�i�v,Ks�n���A#܈R~��"�{�(V�]�[l#	0r맶��э�-�P�T�.d��?��hz`����xQ*yEa��|����5��� xD�`��q���ę�ρ����5���5#2n����ǃa�wI��fk9�Vd� `m��߃�G��A ��X��B���#+�Җ$�O���
 9|ڀ�������o��vM_H���ͭ)̰Ħ���G>R�%���� :.�D|�h�(nwBk ��3�Xy�z^}1�����.۩�$�)�bʱ�A	5}���=�DNd!v>m��K�o-{at���Xe/������4�Q$�����bu��p� ����DP�R=�#?�0�!,#���cd��-N�A
<td.����I4��, L��aRt�ܭ�����3�v�oGb
G
�q��5 ��-U���x�	1��$*�^�B-
N��(o��rU���u�>�n@�wW����!����Μ{��&2O���� �iO�f�%�e`��hD�Az �PU���Ȍl������|�TP��A�{S��w!��_�;aӖ4�ř3W/�&O���u
��0������;
UF2�)��R,��h*��FAZ��w�sl65�����-4s�}���V[P0<�z�Χ���ᙢ� 'k3�n�{,8�d���{���Ey�_\����a��@�*����%�7���FCh��6�
��	�=����8���C�P�)�?�X���/��hF&T��ߠY�̾�^yi�:���*vE�-�d�+��+O����4��4�����>�*j��-#���{�b!Z�ƣDR�Ś4�L�1����G/+
���q���d0���پG`��H-K&���)��d(�ck�gglP�N7�
�@՘�f�C.��V17����0�GV､&���j^c��h���H�һz?Iwa>i�l�S/8����n�$x6�3�!��Ĥp����_��f�%� cB|���a��?�oѕB6� �1kn��5���r��dg��Q|���3�{E�R\NN����,�*�v��$���W4��}�L����e�P��sV�|b�~G2�ξ�H�w�zo�v0MdA/����O��k�@�3�X1w���\S��T�]��N
v���������d��8���tX �r���U�C�s����t���m��ԈI).Զ�;ȆI��$��?`�+����A�����+R{mQ���b-|� �쥤>YK�(m�Sc\H���;(�65>Y��S�B.`�^�UC�R�Ee�1���!�G��r�m��{�4�/�LB3)g���8O�7'ů�76.Q�mt9�%+�`�b�V��T�3�#	3��u������V���/��Ch���A�x2=��n�{��L�]���� l�{1?K/L�x�Իz�գ�R�ꬵ�d���>��v�*L��E&�$.M��0b\�A yjcg�7�6��q���Uvt������Z��WC��,$�d�~����*m����Ȏ�.�U�^�@w@�z�B�;8eG�ש~�Y�0c�NŨJI!k/�0~�%.��Z��R�e�1���UnK���Дc@��`�^�|P���H-����3��A�q�W�*
�j��i��~[��o=���$�b�
&���P.��t~����(�-���-4>h��o����"е�f���ыmPO�)%��L�q�j��lEF[3=��A3sn/����Y��6���l��#^�՞�`V�/v��	s�\!��#���W�nâ˂*�3���C!��v���Z[{P��j�dg4�C��w����
#�,FfjkH7>�*g�*��"'3��U+����Ħ�F�)��dTb�����8�nJ<�L#��8j��>�aA��2X���p0�G�)�Am�|yH� �2+=��T����PUi���)Ei{��s����{Wp6_��R2t�%��ڝy��j�����S��	�n�0����\ ai�8��&7=	"�D�ϑ��B��~�KWv��/"��z���M��²��h:EU|m�-Y4"�X1,�l��Ŀ�*��W:�.�X���l����d.,/��ԭs�p|��O���� ���xL��Ӆɶ�����ۢypr����v`�ݏ0�X�Ϟ 	\ �u
�ȓ��t�)~�;�=un�ʲ7�@�p���U�[��>���Φ���;�5i��y{*H�
�h�T��J��r鼛������y]S���^�B�MV&��E�ZXw�略�I��+��W�-�"e�����Z��+�b�=���Q(��~���n�Ё��Yd2�/���R����	`��d6Lj9T���a��������lF�j��f�p<���I*��Pv�gVz����h6K���"K.�i n����� q�n��a gm�teZ�K�]��P�
���'��Z��'�"a���a~��}���[酂þP��zݷcT4OZDƶ�7�̭��W�]̓is��o��y�n0�4��땲�b�kP�q&� 1���1Q�6�X�?�]g�
��4��:��ؘKx�f�;BBc/�w�X�[O���t�ts���Jt�}��W��
�R|��b>ר0>0�p��X	�Q5R���_|�ȋ��<����C������������UD��j`�m h-nB����ߕ��خ�A��� ��
e��a��Tf*}#+|���|:���"�6O��~�I,g�"f��<w����&jA@$��,ƨ��8�uʹw�f��`vߍK��M~���[Ud�r9Ӣ��猥��j����Ӭfz7/�:=�2�4C,�6��~��D9Rn{���[���q*�-�n}���K�EqDGOX�7���!�� ���.Kƣ(��v��:�<�ů�6��)���NLc���;�OY���U�b�f�K�-�c�xW
�L�aw�j44�D�BZ�,���C �o@C���	�L%r������ʋ��;k�˺�.���&��Z��{R���o�Z������P$���v(�V��q���|��r��w�6����?�.�D�j@����RG�������U#h!���;�uc�����Q��"jd��?g���@hD�֝�b�����ܮ���y�n�C_į�HA�*�pwU��z��A�y�: �*�@�=�Z�mE�@=��?pwS X�}���eF;_���|Q�*���fx�X��0�FX԰6��i�Ƙ#�J��3M�EiM>�5�|�C�ԥ�j[]n!�2�g� �,N8�5��P����<��;ԇ��&S�.�7���k�RlK��xho�R*���v�-U��Eb�5��Y�{2s��F�#�����G�6�g���}��*e��;�A�_��1��3���#������$��=9{��s��<�����5\��O�8�&�D��C+�J�)�3h�/��+����h�t5|�m9�qX�z����Fzqr��K�L�ũ�u�,��D� ��rwy��H���#���3˹$q��} ��鑢��P�_K2+ ����M*���j$��bd|{T+3M�|x_u��C���;ƽO�@_r��\���Kt"�d�(�"<���i�l(�$�F
mh?(BD������ϋl=�M��$,l٣1pCM�������uǟ��;&��S���N�B�+�sQF���un���x�ŷ;h�E{2�#�H�w}����Y¹1%"��ZV�F����uRom�炆,Z�3����������t�%�#�$�!QJ�5k�nNT���I���9���۱�����OIͭ�b�����K��e|9�Ba�%�T1WP{��-P��_I1=� �xH��%/�O���QC�o��1`��JHea
*�(n+����8,��ۡ�l�� p ��"Þ;���g�~�X��Ϲ�o�]N����r��d7��C`G�!I~j����\=⊎��yq����H��iExaB����jķ3������|�c2���a��j�6W�.�.s�A�u ��زf8b[Z�]+5:U��i���\���RW@Z��
_��8z�DӒ����0ǲ��c�r`�M3����G�s���qz�k-RX����:9]+��q=�߀?j8�E����f�8*���'��u����a��o����k7�-z��LЋSN��E���O5��{�D�G\�S��ZpV�;���G� �Ȼ�k<�uB�q4|��>�4��[�;)*�oU�aWO���<��v���@Ǩ��Y��x���#��&[��M�rN}�y���W�5�ʔ�'����Y;��+_�C�Ç�횥�R��p�+Ӡ����ј�b�av+�O҂d�5Y/����t���ɕ��3��dC\B�T�z�ɦl��9[eXi�V��DC?p�&�{�X��w�$�;��%�JY��o댣�̜O^И.*�E�����*�JkV��9��u���*�&^~�៲�ec�Q��2v{� ��s'W�tkI�}��7�;�[��ZN�;�nC�����A�&`t��?��\�_��-;	�>����9�?ȧ�����Π��a�}�جK����޴:���Rڼ���
꿯n�	��FLX��ȚP2��~dʷ�B�t&"z8p^���F��x���)XQ�yl�a���9#i��_��݋mTj��	5l��3W�q�a�'��N�G¨��b���/
m���4�����<���g�G<H�Og��T7�c�,�Z�p�˅��A���x�?6 ��X��n����ם��.]<������0KQt����]h�2�/E�7m/�!d�V^���?52i�$`{���*�x劻�'�^�!�T�Y�ɛ�ns�n�CGa��.�-���1��MZ춿;�S����`������O@���P_w�7 �\��w@�#0�W��"<
�&k��:���IT�����������=f��}p�79|���/��sϜ��%埶J�ښ'�ߢG.�kͳ�g�ԧ3��p�x�c�'�����\���3^[u�8(�kJ����\&9��0{._���Eփe�q���9U�ß�0�ݝq�b���)?p�$3��ǑT�2�=��;?��L�U�=��{e��f����V4!ۚ��|ʅ_:��(@?���Ng"s����N�p$�y���5�Й)Lr�4�|y�\m���\������N�A�������h�{�5;�0r.'�V�����WY��V��1(G�����Gq�fw��z�<E�Wf/.����iT�>7� ��&VGBf�>m��l.���K����©���ظb<�w���3i9"��V>f�3X��;��$~G��CP� ^ݜm&�~�P&������*����!�����_�((�4Bvȼ�'�Us����JYރH�S�U��	:Xc*7&_��36�� �y�s0Bg]�+���hs�g����d�������VXU�B]\��t[P~�*q��^�JpC�Q��ZY�o_��"��6�Y��<�9�܈�>ƽq�������#/h����S������=�4Y�����,KDC`��	tL�ɢ��mP�L�ף�E��7��|����SG���j��ν��9_a����I
Ql�7�
y-V���-�.M6T��&g��Ѫ��:(��S�x@ƨj�d��w��241�`޹�)}4�	�hN��>[�즇�,��$���1>�Ywۜhd�t
^��{�N�_��W�X��<�Ѧ�(Ȉ�&���S���# ��HuB�,���%��`�M�w��T�HN��2GcY�vH�y���uY�����7�$2Ѝ�g�6��#?�Mż��
�#��C�y�'�~�m� �C)k����gL��B��)Y���'� x#������_/��~zW7a�и��ޝz��}3`��W�6�?^�XZz_�V�%TҨx�˱��O4u�g�8E�%2��}f2~��ύ!��N)��q'Y9˞����.O):ќ^^���[�@N���'q��<i��PA������8�!��u�3���M�^k����^��j��u��8���a�z$��� ��x�# S�n +))DEW
���W�ODϯ��o���A�S��U�7�g9a����\��"a�nS���d�1S겝�*PX�װnzFk����Q R����UO����5�g���,�״��{d��z��ùq���Z��{��0l�G����x���5�U1�L�~���.@W�N����NA2"Օ�㯎�Vo���R�sKC����V�c�8s��n+;F씶��	=-����>�g�`'y4�f�Лs,��b��`iBãq��W�|��JW��~��1G����XOd6A�.y� ��J�~UyDeSJkY̗N�Z�o��pe�5�����Qa(�Ԡ��u�&lj���RØ���ǔL�0b�DRX�}�G���ߞ�.�MkS٦$y�Ĩ�5+Iu��G^���Ӭ�)`��C�z���BޢQw�m�;��#�״2z
_V|��v�7a���
����N�-��4E��iGD�A�����B>^�X�^J�*��&����~������j��&ސ������|���RRn���w|���&[�zd8`d�P"V�������Ƚ�0�M#1�녵R�
Y�Yu�)
�%Y�y��'�t�8�Vii֖a��c-3pM�[Z�Q��x�%w�ٶ�T�_.@�l�ۗ��Zmw�;����?DM�t�}U��\O�ۢ�|�2�s̀�����х#҃�u��_�R�Z�#��}�q�N��GE�`���H�o��>$������7��>���+s8����b���r͢�>7�m�o�lȟZTga}���_��Z�0�!pXV����~;���O�M�&����M'u}��+C3�"�T�Ĕ�n��ZM��~^wWvf a��ߚ������@[�Ո1�+�)s��*���T*t�5[Ǵ�2�n�6ϝ/߫XB�U{�W0��y��3`��[fi�Dƛ�l>�d�P����R[�	ϐ�)��Đ���*�^^5���.�Mۋ�=n&xoȳ��1�=l|�k��Dq���E�/B��BG���=���j��m7��d��%��c�l�s]���{�}'Ԃ�f�����]�>��O���s�Mv'�*�� ��5�mN�Hgc8 �|k�AǙ��O^ %9Y�0͠�)��6xx�$;�M?�5��p��.������=ϔ>�I��TP�̳���]���`n�>:m����z+H��Q؋>�0_Q^y�(�gfL�ܰ�@����1e-x���LN>G&�ǽ4���*,�xc彭K�!J�<"�}^O�-��,���8bɾy�����G���p�Ɋ�<��7���9�VZ1��\�����h����j��Pgi���Ƒ�Wjщ�F9`�Q�
��'�,��7���9��{
߲��н�_
׶��,LD�H�wq�sW8��:��8 
��*y��2܋7Y�I}^��(�lK��֨
�A�#3ńV���ϯJ��#Q#J �i��nD�����s�~rw������\e{�[�0H��uA���(�<\����T�K(xQ���4�p JE{�XvÄ�#���&�U@l�W���w�,G���<]���J+�g���]�H��Z�[��r%���
U,a��ѳJUK���/i�G���P݈�1��jll�I��'3@G .�H��wE.O�n�p�ݬnE)���>�O�i���F֧��Ұ>�[�*���f�̪�&���I��5����w�#��Zlņ"��g·�Q�+���Lz'�R/����=�e06���Ϛ��@5X�㺄26� ,�X�{�<ϯ{�ӻE'~�L��FE�g������u��)�$(�Yz�B�5r��ڳ��̕��?"<��z�=f����6�:z�%�M��Z���u�����͡�]�pu�@���}��1Q���d����_�Y� �8{����li��>���ܝ	���-)�
p��[Yn���qn��k3��s|����h6�iY����3	�S�|׻���Y��G��ٵ�6]�2͂��ij�A|���A�:��b�У�<{ľ:�m�B r��<B:+����Q��� K�[JsG)�Ay���.�<W0C�6k8����b���\s� �sot��ېv�ד�N?�Y���6V��9��G)(9�&��4�o�hQ��yE��2�Ԍ$H�#W���Aw���}���mRS��(3��$���u�1���2�%W� C��N�jfi2���yzyۡ�>\;�K�b�Q�iڣ��\�w�@���� ���n�f����]V)���F7��a�$��vB�"aL��L�͟���tL��J�%R���ω$~-�:1̑=���ޒN�_Uz
dW���W����s�>�T�g�W��S?2L{
��*�rZ��B��ʷ%���(k%�m3�j�/���j0�ځ�Ӓ��X,�$M
s0;�C&�B��z��T<�|��,�-r3@�æ�Ax9&��%I^�]Fv���L��'<���.8$�*��D�3�I6�A
��O�t��C<�Ɉ	)kT��猂���ieV�8cw8Q�[A���qY3��k�>�i�Pl�H*'9(oM�����k֎v�I1�/'z��`
4���9��s07�D�.�y0a)��d��=	Ǳ�4�5X⪑�1�[ͥ{+"��ˈ^�N��_�R�((�~�"\�v��S*Ǳ���k河R)��{�DC
�g�8��b
c�iX�׷k7��H�l,C����y������=/!�G�8e�:�9Vn+�k����Od�ݳ��%M2��x�Zq)h��U��ӖT9H$�0#Ƿ��Wq6��J�A��Q��מ��nwKټ�P��
��J�ac}�H���=d-cֵ`S�����p�#�9{( JR�H�V�k�܆�sR;������+�>eI�~"�ɍ�\��˨�U�Y�jٖI�����KB�f�4���:�!D�"G�q4���$��Uժ��O�W���O��n�@����=�-� �AC��U��a�{t��ʘSNM���;	[������}�eoXd�20��fY�X���ty}�|/�2	�D2�J��� cG\|~�E�]��{u��v�a-v�����,z��ڴT���B#�{��=m�ς��/HR�4��q����ts+�#�i��V��>S� -��\}/K���.�i�	�U�ͅ�E荒DB�)V�ꓒ@�������������$h������"8+�{�=ʜ�8{��=��#�J�1Q�v�"KsoA�����g��P��e���H�숾p��K1�,BP�Gta�'��F������+�Ou���鰟�ճv���Ê�TE��I_@�ʺ��f���,�_��ĝ�A��&��t��{�ܠ�W��^�����,L�g�LLi6���S��й��"�K�q��V��}y��yy�F�����^�1����~!l�a�c�k�����s{�m�b�I�F!�⟃ӳBH7e�N.�.�!�sQ�v6�ߋ��y�`"{Q�������lO6���5-,��<V��F��i��:�%�#I�����^���a����(����0�B2���0�N���%�h�:�C*T���m5�c�C���,�vW��A�nh��Sp�~��S�T�bH�a�[����D��ӊO1�z����`������[&�,�;�n����5�Ł�BkN���� i7��^����ɠ򴟢9�}V?&�(zf9�Y��u��ګ��f��Bz*�D3?U(+X���o����T�4�7���[��6�£*�*p/u�#���ːm�8����]$rj������s��e�� "kd�o^����f��>!���\���ɬ-��uv��?	K���}�ln�8@Ҙ͆M�ٿ��0�M�1Y�8t��5���DE���j������8�Q�r~���CL���3��p��̔r���Hx�7�I�_?��l��U�������,`�p4�&�y��3�
���<xӬ�>q5ca�x�d�C��X�I��Vɜ���?3\��ť�9e��%p� !�Sl��ۡ���!�_�ox1;��\A�4�%Ӂ�B ^,�C��T��AM��3T9��������;�F���)2ڿ�\�<�8LL|�����p"Q/f3��ؚir��Yբ,�`��P���*áj��f�BX{;�x�T�kqhvK^�&Z*��߁Ɯ�Ú��'B}�v�
�h�H�B�,�uǠ��|��K,«JFz��O���M#"�P����8b��<DkR�s8V�2�M�V�@�3���[o[m���ЎG�����GD;:Ҫ�X�-�o^],EYS9�'�8�Z�ؼ��k"p�;/^5�r �V>�T������i�D��SI�W���s$tB�ƘO!�/y伔������FLņ�T����+�W`kh�t'wG:�SZ6l�۷�8t�EG}�]B�>
qe4�@���n.J@]^쫌ɓ�e����u
�Zێ��;g�����I�V�H(�| р�c1z�"K�b>]���M�8q��L�������f�� w;�����$,tc�������a�8ğ���t��cJ�˥	Ñ�IM;��`�/�!�1sZR���j�*`���Cp�J	���G"��z��8��~���.a�$�:�<�DH��Wǐu$��>��R�J)M�҅a[��eU���ٯ~=4pI���# ��/*K�?mR�j��.�;�D��d���R9Imçſ�.�`/p����.�2�'J�����v��$�Q�߽P��D?�qP46_� ���e<�>�b���	�h⫣��W��r>π���'�S� ��T��\�����"�|r\�r6�ا\�>�M�Ȅ�>�m�E_�y��9�	���.� t�5d�n^gm)���8�C�8���$NE%~���u��d�=�P��<���/�\x�=��6�B�2D�K�0��c���;'���N]������0�(O�1A����5�;Qw�5z�����D9�)Z6lE a����=�_���O$L؀.���{�kAȵ\FƮd�E����h��M�H���18+��7V70��g�D<�uA��!�le�.o�M�sDMy�6��!ʫ2l��4���m��8�d��#�l+�`d�V6��y]���I�3fR#���[�]������T���b7\����~��$g]��6҇�����IܪS(�B���	�����l��,A���֫���ʩk`��%C���{8�<)���{q-�zZA��W�e�*�xܴ����֖d:s�(������OT�bl�Sx�nf�Gc�ڝӮ�P�>���݊��jTM�sG���s��Z��m�(����*�\����6��ʓx}T/�U�@#F�R�6]-�Q�CU�.��2k%:��m�H���{�?aK�D�Vs�bw���e!T�n!�giȰѬG�X����̵?�zdEA��V���4��=*K�Uw��\���+�Y�d�5��}�y�� ���䷨����&�^��liz)4 �V�q%�9�����^��A
s����G:�·?N!��;6�L���z��>�ȼym~�Ă���U�аLR;̎ve���^���_]=G��n�D(��8�/u��z�ևJq��9�}i����Y�䖼�tD�T]h����+�h�	dU�� ���@��u�� ��P�_=j�*�n�\�c���˫�|��&��5(ˈ�����X�{"5�)���غ�*�9������'1�苂�@VV��EҲW~�l�
�v��H��R���(�s�`J(�}�=Z�x9����w���6#��������
2�"I]�_����OL���a��܏�̷���[�L�F7,U[hmJ6�Ff؝1�����Aט��0|����h�W$�N�*|`�8�l*��N���"h�~AoD`�cR��9g�B<�\��g-�A!��<[K#24�3�ު�-Ą-}C���9@�J~,�7�d:u�����5P�mw�;)�x��H���bZb��/��g\r�cɃ�΀6�جfA_��(x^���;��N7����
M�-�N�$D�^J�R������l�$�3�Pd������_�hk�b�j��y>�t1�N��K��lI��2��=��A{ѭYR�/�I+of<<�M��}9�#��
�H2���"��_N7�9�<d�Rb+�alL���.#�o&Hytx"�m+���,0c�럡X�BΫ��V����c�R��!cv]�]ܯV-�W����Y��P�c�. ��,���ϥ[e p&�K.c�f�&���SV���c�|�k2����@���ۭ[]���[�����!G���������P@���M9������ޝ�����'8ֈ��Zff��7�������T����^��ur�:l�M+�*Э[x�b{�^�˵����O@�U���'��i��%��)�k�B��_"RԹ���>b%�b��xe��a[|Z�{�FI�C9�4"}����8�P��U'���RT(=6{�������!�*�ſ�Q�QK1I\M���g��y��f��Yr��w0��5�#���Q�cvO$�Tqx ;s��v<� '�Wi�-�cs��wF�egoZR~<þ�������w6#Z���e��ɛ�j�E�fe� �I̛t	���IS�cD'�$�"ʦ�dMg$_��H����Ht�q��,���g�RN'-�Zn�r�Ǎ5�l�~�f�W���=|�.�I��K��w�u��JaS�`�6��MIP�ǃE��|7+�=������$A�⏨�!������.��m���ܚa��c��G~w�]���'-HVp�pm���}�!x�3�����4��(��J�Te{�`�6��ք,����Ӊ�I�~����Hz�8-q����}nI�j҈�Jާ)����`y@�D�6�����c'	�[
��[ZH�X�m:�z��o&P�X[?�d`3�݄�Q	����n���S%(�M����B?��C�5�7�,����ɍ��Y/��`)�ri{}�G���^���C�D�� DK�]�+��L���2�ī��f�㤏{��P����-d�Lh�׋�>o��rqbք�3T~�}H���]�yO~�N� �~ni��S�݋�@559�b��n�����21�/����I��zYB?fP�:��l*t�%]&ut�Nq�U��x��mخp(�	[T�s�g��X���A����;��l{����- �q#C[!�C����K�����{q�n9[^r�az��B�#��_�q��2cjH���χ���k���0E�ձ&��a���izԅ|�d�@������p�����B8�?�Q��e{!��#�&��,��bP�v��Sa���×����i ��q�����W����
�:f	5�����o�Q��Zl�Rޮ��z���o�0�w�G��鴋�K�H��2"3�7���e/d�'�--�-�1cb¥�o{����{#��>�3ƪ.�4�NK����a�-�+�1�e4��gC��4cz4�n�:w8�9�|`�|����-ޏ ~Pn���>}�c��&Ò#�o�	��2�Ė���L��C:��i��/����F5��y���?dm)�*l�2�p[�}-^���@<U�(Ɇ�K�k�r���`1�%L�7v��yE)���n��t�q��3#�]k1��b+e������`b4�����[���m~��Ի�k�4X�aZc�M���v�������0���Ͽs�1�5}���rmS`.)�u�����Qnk����I>�����X�m�Fy�A5�
�Y��7xڍ~����x}��B�0RᨄL�Ώ��7��p���
��k-�Y��>W�Ӌ,_Щht���b���}7��5ܾ�q��(���M�����^�fG�e�R�JV����2��J�g��X?@'�ٜL�9qp �#NX��x��W�����02ޟ���{����a�H�Q����⢅��F8��x��۳��>_�׭7\�8���
��Bޚ����A9�;к�F'��94Ҁk��I[��ԟ�q0�{N�"/�#:����T���}�YB��jn.wes�IQ`z�
�h�%@�Su.���#��<M���1DƂt-2�������~[*~tJ���.�����N{%��ճ��E��h2(-/�>�Pv���K8����d+w�n(Ջ�o�;	�Ln�&�E��:�[��s�#�nW�y��}M�jʛ���D���=ƽ^�N-nO����
����z~�b"hQKE�Ro+��Z�jE���A����Mz��;���#��y��plN�Y���Х,|=��߯�v��#jC��*Tx�g����VrP��25j28�p�%�S�뷐2�e���d�'Q�б��V �иh�FĹhj���;O ̡1���mwSQ%�Q���E*ʹ���u|34��o+UX"0z� �}я�}�K�	�(`{:�(�u/�	س�����:+�ݐ!��c�&���A�D��'92j��L�Gx�
���̟��_��碂�~��G�~0V�P4U$ğ��ڑ� ����}��J�^k��!t�Q��e��r2�i�P�(��r��Ts��Z*%�W@��Ԁ0�J��%�͵nu��>m����`�n�s0v��˺�ƴ��?h��� 2��t\���)O���Ũ=Χ&?��59����zAl�&�oth�%f@d�q�CQ�[�ۦ_��J��w7����S�����������)� G���3�v���؞���۬�,!��_Q�<��u�w��xP���N�a �,ķ��+��&�p܎�X��p�%`|�Qx�~�r����*�49��w��b�h����-]/M���m+�Ȓi�j(�W sd�/�T��^/�䒊����h�� �^\�i뗶��׊���Z(�����0K�A}$@��$����N�:[pst��i(dmV(��`��t�DD�&w��3)˗ ��DĞ�}�G�xh%��Z�`[{�Y��h t�.���.����H���Ϛ̲���v��FEO���hn�-|�!멩IO�EY�ӌN�3+&6��UR��J��ğ�-��u�̍�@���oH��]|MI_�%�3K�l��ʍ N�\��y.�	��,�z����� L��(�v~�$�c^#���g��H��������o��hI���xo�bd��1
/k#��T8\���9<8*X�y����P+������˓z����
�=[>���� �Y���_��6��`��3��$�o�o�GvY�&�hP�����7"��j�.�Uִ #