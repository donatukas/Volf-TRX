��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.yu�=�6B����刮��>��h���!�2J�X��BC�P��4jgLip"ח��ކ2�%ؑtG���?�H3�o/G݉�ɟ�x7�D��T1F��HkH��+����ԏk�2�h{l�?�E�x?��*�%�V��x-}G��BBf�ee}�]��AuTX��x 8O�2��,5� �$��8{�C"(w!���.�g�����MT�%v@�r6�۷��� ����sM��Z��3HI%��I����$}��hp.�7��������
�g���5�QE��*���R����s�Aͦ�o�IJ#�(m�B�ߖ�)�v�>�̥��p�bxau�d#��&i�h���U �ve��/�)x����j�l��oB��@M��uMIĳy�A3��+�{��O�&G�;g��B����KP�Ŋ��n�]I>�� 21&�f��h��	I9`&�F�$}rs�J&�~����i^���mni��fJ���|�G�|U�w������@�/"�AK_���
��G�A]Bd��@��B,�x�5|����R4P���!# �����n�ޣ���>Xdf1�y�&���ma�GH~�b��L��@yi�g��$S�T?+�*���n)� #��U���Gh�/V�*9�!��i1��h�?i*��Y�KjM|�PT�i�y;��kί��j��o�/��+�m��K"�[M���������zà�gq;o����.�8��I8�]�Rg=�=�C׺���(����{=���	;�R�]M�>cF�ru	��õ|�pX����[P9�?>�l�#�'V8���>�9Kv�<���7�E#�s�\����a�L�ۉ��d1�5�{�u��y��ʇ��ͺ�a]/�S=G=BO��4V����$��Nm�������W ��.xp�!�)}��`�{l��aQ�Rtc��$q���گ��)�)JS���؄��!R���8��f�ங�.�1��ts3������ ��*�\���u���0b�#��1.XU7�����C<���4�dZVX?P?G��M(�w�)���'7!|x�������40��Q�M�������ϖE�`��I��dV��yz�M��q�� �8��w_÷:'h�r�����V�.r�lf�Y�{2ا���g��K�R4��o?��$�~'k�v"%02�����<޸�D�O��@�� ��І��_���������@��� �����P
�F���Jӝ��/N����!�Q�U�D��A�ц
���Z��� D:�&����$נc���㲙�kze+c,E��o��2|�Ho �^/㼬[i%�)��$R�R:�6F����5 ���$.ʟ�o=�ն{�>�87�� ���	�#�����m{���p>�W��<��B�|!ŵ?Ï��`�p[���)t�脧�R;g$S�	�h�Pg�Q�Lu+^m6����Rh�3��g@e��@`a�Au����"�u���c��@����/��m�b�t�c6�0\r��b����dK	sP
"��q�V�q�f�a`D��%O!��)���E��c���b�M
��(�⍮���B�C�+h~X��kN$�
d|�f�����թ�m<�S{��E�F��MTS��X��]�@ �{Q�'q�S�gXSt`�h_���Z�Ic���|	А���eD�y{eG�T�9���,�������	���ٚ�����"�� K����\��+ycA��<9S��-�C��f>k^j@�@����B7C�ޚ�����7���hVGEc3_���=�'v����{ H��.��WO��kX��v4V���a�"Kԅ��'8S�6��mp?6��O�fk�t�c���\��l4������|��	�N,i�a�Z��]���W��&K�7rz��{Dy�;�u��	��Y���C�Y�nt��1צlxQ����ߤR���in��k��EV�}��%�	3,ط+�,dZ��y�A��Ѡ�otg�!��\�`��$>v@�m.�[��:b9{�o82��+y�C��m���Ј>�i�a,��ch���{&77�'�;4Z�"���C`���UbP`nW|��:n�;|u���f��O�e<+���~���RX�|�������h�i٬�/�,�5v���"= 2���AM�B�]U�'�7-y�Kb�PAr��UȴM�������!HX+�5��\���s'3����w�򩅑��&��ǧ�)긋�r�aP���7~;�U�e���+��ѷ�L~�~z�{F�'
�Π\����Ƽ������>��yɗ^R���v��g0$����*��`�%)�1��͑��J��yӫ`X���
��r��ˈ�Rx����A`�[%�5�$,���%�׆;�. ��C�~s��]�����Sq ��kv6-��|Q�Jb["5�5�8\��~7"���F�KӞ�|=kAz���r�X�C�o�;�l���W��px|��o��(�kn�k>��;N�M�f�͌����H��Ig2y�7U�U����
�u�b5-�Xzi��z騊z�"��<����e�����|�yB�z�:AH��37;����+7_�@M�ew��B-c`�ڂ�U�=;
W����/Ȼ�d�7�I���BV��upu����/87����{��Wp��BB,R� T	�_�76����j�������é(�PհT�U��|:�Hz���!W+v�5�E�$�H�lw�-�j �K�S����m{�es
��E�A��k|ֵ�`=��FVu��w��cb����{���_nU9&�ʷ�����?9�E�R���?e�?���X{��ff��潶�:�L�dF���%��Lr�C����� �}2���Ӻ>��D!��m��Vtsz��2U�(���x�c����{nS�j���}����0�ϲc��b/#0�?W�@��iU��Y�l���<�g|�Y�}�D�\�:��z(��j�eOTyܐ��E�YQ���:�O�kV-$�UuRP�<t\������Cb��w�u��*���|RW����a��I?0cC"m#F9�,���	����{�Aݎ�1g�0��r�~�����}�8��*I�t�ŋ����qs8*A��R ��Lka��T��0o��ǯ�<�þR�;�хC.gv=��L#@K����#�/�0����
��;��Y�~� J���5�Ӑ�´�k�i�{��a��hy�Oc���'z��=&?ԅ�i���M�B��K��se����bUW�ڰ�r٠x$����Ś$�����;�9����/���\���!��֜��Ɓz�:��}���p�Y1��	��( G*<8�׋%Ϊ�z�i��&�%��;���zvY�Z魋G�t���P�OPU�t:�} ��KQ¨t�����GF��R��Y�^M���3Y2��@��-�U,FlF�42kf���ES��r5h�D��T�nKk͒|����m�6�UĆ(V�7�{����ϸ������7��P�sp�K#��Am�����y	����٦Z�<d���U��iFz�� *�Vk,�+]��w�_ Z^��4_��+���IѼ1�k��V��	�[z�B���g#�e(���DlYv2���{\���3e]�U��V@U��wHP��RS���~�A�Wb$�-�����FzA�~�T�j�c���� ��u8���쇒�6�o���]A9��O>��A�̒���z���h'5A�"��X�bߜ���M#�EZ�3s- ��"$]_�{ß�^�L�H �if ��ig���f�̮!���)^~:�F��o�]v�xpz��}|�V��|�-�Qn{d7z�����2�Td���a������T{%;�p��u��&%��3�t�3�Ei/���>',��ٗ�G�C'h0�M8qHq�s���l�N�O&Z)Ϥ�*c�RX��B'}Gշe��e��E噻�먋^�F	3�ܤ��;�Y�u���5�����9�7t��!�~��1�e�ˡ�[����5_� ��݉�G߀������3�t���Q��F@�uDr��{��t�ٽ�$&�i�
%�5 g�V���ȶ��t�k͈�p�`��Tya��>�sq+a�3��i����?Av����u�Z�|��<��]�'�c5C�`t����:�Ir7�5�m[�*e�p�#Q<!�1,��`xẙm���9�8�6�c7䩜�CϜ|"#���G}�g����b�NVhÓ�� �� +��m��B�U�T�턠1]�P��4�'����#	h��3h0_�-�ҩ�U��Z����1u���F�uUgo��i���pG ^�CxD�*�Y8�V����6���}��M!�8Wy�N��p�'����F�f��p��L��mը+)\q,�{��[���gɺ��lzl�>b�h�IH.�L�kqM4Ke�(w����_)R���NI�c��1;;�t#�G|?h:�m��*e�WMr�ԝ�2Z�s/�P
���Iݴ腠��e`^���ٺ��7Cx-]O��u�o�#أ_�l����YM�>��(+i�}⏕���K|��8"Ċ�ٖP�Yݦ�=���&�ߥ'0A�b�0�V!R�LT(0���G���_Q(}��/�W,�Y�є�[gp{p#tƅ�F�f$~b�z��ߘb:x�:=5>��jq*Z���7q��( ���;KM7����w�v�>� ��R���$!�&KCb��Q+�~wY��J�o�|A��o�PLNk5�=�
�\�UU�6`y�{�=�'f,�BIw�/Z��8X�I�����D``�{ឆ8�l�C�f6շ^R==sD�A3F�4e��<-!]�R	V�I�1!����@١J+�P���M�_���[�!;�DTE��{ 8�\}��:[�-����i�Ѝ��AA�UG�"S�9�3љ߂���T���2�hj�v��֏p�ζN3�M׈n)������6;7�3[��!l�UA`^p6��Q�U�8�&	���[�Dj+g:ↀ	�S�C7���4*�:	&�^\��ӄ��7nC�f��/�ʬ<��-�,b��4�����:���n�W��q�x���M�!y

��3y������6�a�*��GN���)��V���(Mi�� NH���W�rd�9K�TS.�ziLC�WD�G[6�}�40�yB�׺G��#
z)�-9L���D��^ؠ|��ݫ�k�1�m�˵U` �B����D��ۮ��@
����i��xY�)<2qk�	�Ѕ8U��x�I�[󷸩VD�6K��"����x�'��^�(5h��Ԗ="��b)0����}�F�.�=H��@�Qݒ���U�\<!D��&Bko�SF��.�芜ԮDE?�� Y?��dN���ʙ�Q_"PJ��)��y�uKW�3E���WC�{�w�i�a�a�''*�����F�6�Pf�dO}d����M��j��>C7�"e���{;�ԋ�z=L9�p�zH%ߠǧܿ@-h����r��{��BA���6H!g��;)�W��c
a�c��b<�<���%o#)��0�G�xd�v݈Q�Мόסw�a<�.G���[����W:��1����_?D)�rd��S ��4� �,j6l�*Y4��s�i�
���ҳ~�_�$@����I˲[��-���AF�W�����n�WXO�Xr!`L���I&U�z.��qT�C�I��\���K=��?{��H���B�4`<~wdw�"�C̊J	�9�+ʽf�4k	3:�2Z(�f0�9��l���lA���(����T���2��H�����U)�-:Ԙjub���}�d��-Zǭ��m��C�4�Mh� ���O9-�_ޥ�yAy�j̓�m�G��x<�|�̴��f�)��N)�HZ�vǍ��u��A_B�%�����V�����TjO��t,��
v�~]
��|�����=NL�d�}C��д,��l����5;�?�NV��y>":� �U�^yo����^I�R-��J��!�k���c����5O�4����~���q�8�4j�y�@�}[I��Q���2�l�8`ᠦ�D�VI9��J[/�N_6���Rd�rw&��,G�|���/@�>��ӯ��W�t�c��bq��C��(��LʺN�~v���*�%C^����N��M��H�N�d�_^����56�B�P�z�A� J�}&!�0@�;��峵	��q���L!��E3�+�Yk��K�Y�>�nwn��?�Y�r�'�I	��O�ؕ�q˻�v�tz:�SsCq!���l�~,AT�P��`�W�7�/�lW���Np'�0���<�S�]�4�#<�l��E�߅�$���	�������_/��ފ	/*2��@V�L��䫈��q{{'RĈKю���5�k���^�rEH�tv	a([�^��a�7k��հ��%G����.#D^L��fz�j)���d���"O�O*��)�6�
���"<���G9�Y�]���pH�\9����7�gK}��H����N�>za�e�ǘ�ƕ�����mo�>]*RMnzM�w=6���)�z��b��ɵh�����$^���~�ћ��wt�!��?L��f[j��~mҖ��i5�+��Y�a��n�S�JQY[�6�tw���+�;�&�5���4���37�W��P
��D��_9����1������`+;���� ng��䲿<��i�'�*n1
�R�~����ᕶxoXW"Sw�ѽ��RV��*���13OB%(�T�������Iᦍ
t`���<��~$e^x!�����J��h�p�e��;?��8D���Q���.�\\�^�'3����-�"쀊��17�FX ��ߵ'7�q:'���A�+�?���m�����Tw`6N(������:�Vzn�r�k�plB��9��Y��3����b]�B���������l�/��0��	I%�E<�=��;hX��[_[��x�Q�`K�l=���x��,�%T0n.�N�e+�ڴ�@9�8�힕�̱!֏�v:�Lp����RV�R��_��[�נ)_�z����n�.�/���P�7�K+o�����U�:��tR761�i�9d-�gQU��欄�P�c���j�0��1��W�m����@��^����G�x�C��ҋZ�����/�`=��a�k�ހ7&�� �NSB�����?m��*):��_��w��z�V%1<Bu<5��p�Ҕ�|x�&�(�wM�b<��ĵ?�T���m�*/�s���I�aL�+�w���c3���b�j�&]Ǘ\)���E�KFf���c맭M�MC����˭6�H�n�t-�N�D$Șc�����v���=�̷�f2�=+i0m&��(n�Dzt��mg��o�]�#���!JN�E}���G�ɣ])����ۼ��!��=�6��vD>�YN �Ϛ
RY��Tq��?����$[z��MK!��)��t 4�\U&G�N?�;�߶�)V�� �������~�AZ���g\��Y(-�����Ih�-�����{�<W��o�j�a� \��(�z<<r�U' �kf�q;���
�G�g�Ӫ>d��-#S#3��z}Q�}Z��A�lCH���v���E�k�<럞�W�x[���{Á~8��|��
Q�d`��-�������w��i��~����0x-g2�:����$�{W���i�M���pɰO���4��8M�/�׫x����ym���+�"�iK^;��^+ߣ�or��+�m��ꘔ�
�˙�S-�-@��\�ʶX8��n\�9��k�t�S�˱�yT4X�s.H��!�a���6W��sk�f�	⧏7G���� �<� (�G۳<�����i������,��죞����7���:�Ut� L�l�̠s�!�.@ ����&��gO��N�u��o�X��r���[	m�¯(H�A��[e�Pp�]:>!��Lf:Oi�w�{�%]�c� ���m�F<n!�[�9���V	|�>�PiF\+��bB2!�"S�f�z��e�0�6����{G�we��R�bk�& 
u=񔰍vZp_r���������oQ��Xb.}�<�^w�Ե�`�������r��X�L�p�	B>i=ivCF����<Jp �C@DW�0�����G�D�K֗TݮC���1��ܾŇ}�8~�HUխ�u�G���;���QAd:�.��U0�C�!�$�Ƒl�cN�|#Z�Ad,ݩ��j���8Jgث�ok��z��/J��1���*���_\�p�e>Dr蹎?A�J�~���Q�j�V�m\�z�17���"�z'�M��?p��X�7ݯԧ�sS-�#�Kgp��Q�Y,��"1ΫH�zUvӌz�B� |+�O�k���yo�#�{ =Z�+9��K������7��ve�y�!@l�QG��y���D�^ �r $�|��zE������ {	�����e�[�#^���jlf��
/U�u�+���@z��.
�������+�w3���(}�j��{V�k2Ʋ�*��W`��y��*���&�����16o��`���|�s��G�T���&U���	&�Mt^��0��s���z^We��N2�s �˂d�*3�O�׌���!�p�����ܻ��pc�:RH�%�.̸[�^���p�&g؟���Ӄ�jۖ�����#Dë��.���UkE`�e�/�۞�?�<0�o6O���F.�b�q�p�A&����]Y���@n8s�V'8	��	�oy��>-ۯ׳�1��ô|��u�f���ߟ����|�<t7_)]�NjuLx:�J4�"<·�酢�W�Ԥ��������y�{��8��c��7S����e�\�����!��F���	�|������m1��!tYFR6xo��Z@3VR�lm�<��.����Spawl��������X�ș^3I����&�q�U��,Zر`���L� �꧁	���m��N�)�Or$�C	C9�M�EY�"���F�h$2{�zk��Y8c���&��4�j�f5X��h� P(]޳�[��3��8���挾�@�Pc]�H��ק`�C-Ֆ���@�/!��G<�P�b�ǽЪA��/�1��H4t
���,�ƒ�����X�>7Z�e��%���Ƙ����zɈ~��s�_������W�"t� t����ӧ>��g/?W{Nr	� c��ݨ��8g��ʗ��I�u^fw���5�jh�5g��cI9�y�J�U��Mç�����X�\�W��H��"�p���+�ᄪ�֌����+xt� (�ac�z�0���9��z���* �r�Ԯ�����Qj#���h��m+R���у�� 'ǃ6�)\���tq>�������5�.來eG�2guVo�'7�t���L�++#(�2k,�:��p4�7m�I�W�!��qN�$zQ�Q�dZ��e?d3F��0�-6��IB� �?��Ky7�%U������GG�������9���CP�@��K�+��逢$f�zJ�5;�*��������\��(���Nf��Ӊ;����p�i�~<\	u�y����yu�����2}��=p�9�?/�d���h���;4q�^ܪ�4Hk"��&��g|{�i^�߮�/�� /���!"������L$�!��I7RY�+�skb��e�N�B�j�Wp޷�P�y�� �z�Ec��fz���m��HWQ���<���7l�]����O��ݟ�e�V����G#��*�B�ԁ��!X����Z�ynU,D�Э�2��7�?Ԫkb��~)�]İ"��l�_}���������m�����Sc~=ɰ�?�����ѧ]ɝʠ=8+�{La�S����!�0�cmx>��X�gʞl�݌�0��	ӁJ&<Z�L���������^�A�	��$�1��*v���
�`n|�� ��=��D�5�FU�tGK=͏����GX�1SDR�oQ�a�����xe�3Э��'p02��9Yh�������!��.���u��t_�-NJ�-W�+ek�e`<�
MX�m���$u���.G9���6՛9cdB?
�=��|fY7�,���r���I��)���hD�6��;��rm�Ɂ�f&�D���9������aW��{6�9����b��Fd��S �.����: h�W�o7�tf�x�4��]�U!�Xm����:������M�B��Xn�}�n�u{�����	_�9�5�@�}[�A���R�5K�y6[���G�!Yu�]�/u����{t(�^Qv��奇1s������+��F5�J���D�ۺ�eDk5�֣{Aqn��F\����f&i��+��npi�h�h�4�a�2c��UV���:�(X�vQk���Tj{��D�uP�6�H����(}Ne`
#Ӭ	��j���������b7��Dѕ7�Ӭ�֮JyZǡ�w�"�h�N\�
�C�P %�-���5�
���#܅�e�j?�+ᄸ&�bz���'{�2D��$5���{ඓK�xX�j_56r`H�c43������I�Ʒh����[�R�9�
��f����v�_7�}��w-�p,hB5�Wl&�Ӂ1}L�wwP��A:�,���f��s&j�`qG�k@�ͬ�]�"�i��#�p`�!�=�oJ��[�h���0��,�� ���I�݃� �z��nB�M�}��.�?�<K�%}��+����ٷE*�3x�3�abuV��~����6ưĢ�8^���CbZ��ZuTV����"�K;�FW��=��|��r�
yZ��K����K9��y��w/������i'˶�b��~��8T�&)�d�e�w����� �g�������>����")m]�y�r���{� J��%�hz*0�8i�8J=$�ę�#�7gs���yN����3��xt�2�}+ث�F�)s�M�q��H�@�Fxq�RS�:E�ر�b%S�E��;�;h��ݳ���ό��|���?s�j�,z���_�����~�[�,jE�b�I�Q��(�='t�i"r���\c�U~̤v��~>fn��D > �1��r�;��%��Պ���3ݧ�KA�9,4��V'ՖEP7N�%��[�ć�����,� !P5S�\o����|�{q�(=�.!�� ��8B�_��1)I�QC��_ӣ	;}?��>�.H��O�C����7��9��_���z:P�4ׄt,�Wd��ba!:���gO<�9����֨�����`g(���2�݃7+k�����9�;��5]�"�<��#�T�j��[�0_��FD"!�V�A�b�X'i�'�B�փ�2��[��'Μ�T��E�N�;]y�)�~�d�۶i�t���,�h���_��{��- ��k̜`zӳm�֣L &��>ؓ��6�O �����w�!�R�w���6q[���#�m�a4��R:�>�}oG凛m� ���+�޻�4��"
��c;�&�>�y*밒:=k�Ȗ��K��E����hk�EU���"�ͨ�6y�t8�G��
��]����1��}&0#M��Qe�`�����c�"��,���q���<\��+�,_7P�%�82�����9�5�E�⢎s��p �<D��Ue>,8Lv�a��?=]u����� ��B�WSRg<�qv������y�R��V��M$��'�I2���F���R{6.�������@SUi�`~*�p&��h���9�S~�{���n�B�dߕ�к��ɤl��Xیq�Ѝ�2}�A8S���S��y��!���,���"�m��qݒ��~�0x�3N��{.(G��	|����j���'�B�s|�х�<��8���ǰ�8EX���0>~��P����Fa��ｘ�ÿ������59�D�©�_��<��h���
(�C�Jk�3	_�@��(��gȌ��T�M�I�x��`q��nKy�^�:u�����������A!/�.��y�4�e솀X'�_QE���l�_�4�p&�8��NFiw�O����jW�qШ�H~���a�|ǀ��|���s��"e�Y	_�5U��8n� !�bU�Cez�9�6��eK��'�]�Y$hC@|0gN��xH��8 ���ׂ�J���� ֭��ni��up�)K�=AX�{�n�	G�N�3}��Km?�cRk�ďj�ܞ�Z��I�s���,��<�x��':���:�)��̍��C��zRAk�i��A�����I����������'�PY�̖��y�6�F��D�P���,�RJP�xE8b��p �Z�<ORɝ�}7��ά�z��r���%yd�/�ak��a#52��&aH�o�\e���/��uG�&�B����D�:��j؟)߷g�Q���5X`%�	�)��L�;kҕ���{K�1}�H_r�Kf�%Gq/��d��u����t�