
module DEBUG2 (
	probe);	

	input	[0:0]	probe;
endmodule
