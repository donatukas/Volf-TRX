��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.��Q�"Gx��F���C9y����.�����i�?eJ�ֶ_v��X��hq.�3(�}� ��,!��a�.K5��FAmK/7 x��թ3>�ڞ23o�{�`�§M�Q���]��j5�֑���8�������9��y����JV��>H���&iU�s~��-��{	�;��[h��`8��%���D��SV֗�ٗd�����*�$k�����Z��'XF:v��2,l���Z��n�����I��ID�j[{�S�Q#Kě�<����&�����
�p�CZ�E����1�/M�[�|؉��u�.g���WJe��%��؛�^}	��_	�	�/��
�)f��;��c�ɇK�j��a�L[A���J�����5T��Ϳ[ۂrr���V$f���C���%s�{�<;���]�f���sC�p=�K@����i�p��^��E�iT[��RNx��BN�ז�-�>,>����2�.|�G���f*2�ך��R���<�o�l�é���A%I���iJ�[�.�h��E�KuR?�g�մm�&.����v�c뤌º� �G�aZXl��Z�X@7����x��f�z�6z\�����w=^�����9M��1��pU˴�����o]�L21��E%�5juK�65�.猣��?�%�y�'�X���~�g�>zv�3�9���-�\�ɥA��sg��x��>����½8��'?`��KY(\��u%�$���CH�Mv�f�=	��x�F��]�5��:��;p{ό�����/Z;8P��f;��������AX��k�\0G��Dd��I�9�o�>E�4��}������%���~qmw�%=�0$i�;�C�P����n�I�r�ͨ���>b�֧�pa5�EQ�k�Mfc��bR��Nf�0E�u��XC���f�L"�P�?�w�;67CJz>��"�u{t��V��!=ɗ\��A����2�9F��~���� IbF��\RgQU<�e��g���=�.a"�H����`�_d5�����b��������^��t��pƆ�'�_�:M���[)(�����]>"��h50�l�D�*�?�}�5��sf����;'����b�	$��uj/u�D������Q;{�����=�<f0���}��ls����n�Ȱ;��?�N�ת]�t��[��	�+zL�A��y*���#���߄1�N��c���3!.�οҝ}8KV>����᫈�i����ǉ_{���@�s����Ѓe=P�n���۔"�]���c:���`q� �t�5���K L�LTT�r��\��f5�U�^z��n�/8�GgS3����9fb&������/�.�z������ON�ɚ�>����B|0�^N��I�4�Ɵ=V��V+ˀ�&@�k�B��$�����=�`I��
��0;�BOQ����S���P�}�S�Wg�I��T�8�X�f��f(:�U�,��9~;�;�V�1��u/s�"��~3I��1�= 
����7PGpQ�U�N�G�{z6�U#�z�9��x浢������-V�P�Pr�;�fQ������#��C��0�:�ޗx��;Wi%��Ӡ|%��
ХX0�K��uCj�~��9��6Ζ����`���5��ZF�G��+]L��*0�#�����(�۔��R����ܧs$��aپ�5Š��M0
(�lȫ������oF#D=�\GE��	�l�;�+�2�7r��!��/���F��s��G�F9U
2����%Q=�C�-)yKٍ��IrQiSi�rU���:�~�.�B�M3�ϖa>C$��6��X���>�cd�\��Q��*N/R@"�0����Ҫ-��
�;z����V�=r�Χ��0���+��n�؉9
�Z[��R��K�f#w^��a�Ĭ�x�֦r��������㱽J��D�Z���LoW���\�ͬ�|M� �b(7�V�CL����e$R��n|����ͪ��_����q�����"�tq�)�,�PN/��d��P