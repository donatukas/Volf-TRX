��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~�f�?|�ў.mh� M_�>/��zTg��P��Y�@��+����t����m"�Q�e���VW=I��K�'�n]�	5���	a>PZ�I¥��Ԑ0���^��r�s��)uD��>˯tp˲O9�U�%���h�#$�Ɯ���Ua��+��cO�p<[�������`=�eH;y��,K�]�#b>�6���Y�з����M �%�R��P��dC��}��(��ܐD$�_��
S-�&oV+DeX���LՓ5F}ƿ�(#��s�eT骀��k��g-��
�4��s�H��G��^y�#C����q�7��]��K��Ӂ ~�C܃���AW���i�u�B=Qw��Jx�I��BKy/�1���� `֩�����b�h�������1��;y����^���Gs�q7V X��P�
��A���:Rfv�C\3CY�Nb�0YXV���:,�>���u����\j��35���^�٧\��߭N�En>��TJ�3���[�L�S�iκ�.�A�R�j*V�E������!�]Z��A�lś���el��K��d��j|SS� �2��/�H㋒�RV�[�O��o��GM���C��(�4�V,#Ɩ��@t\��WH�ړǅ�/�H��D̅q�����uA.:��6՞��$�A7f� �8,t����M,ߵ��c=�%)6_KΝ�=������m��8��;��I����R�}T�o!pT������IHZ��d��u�.��#?k� B�%FE]N{s@9�'���W�ݞ�k�OB��&06�vi�jcr�%��1�X��-�5�<K����SO5סI-��p�n�Op��-�d\��pit��?��9�y��C..�g�Y<F�w���4��	��9����b9=�D@y3�sy����ʻ^�G�@���ii��y��=+�5U��1���Y����I� �u`��M�<�9;1�iA�5��®�%��F��2�	���^���7J�%��(d
mp�Sj[�!�O��_��pL�������$$�Ϣ�3��f&��I'9Ql!��)I0��� ��N��j��U|>s����`�+wgB/��(�r�L��?�M˾�,��h��3Q�כ����������1N3��[yn�z�7D?bzFX�.࡮L.�%"�u|豺wL����MI�*�G�G�1�j�C$�%���g�M���;��Цu��o�����j�v��+����36Y�c�ϙF,�)��^m��N�/3Ӝ����}H=�Yjd�(��R5���{J�@��KK�Ȍ}w9��Y?x--�|=����M�2�F̌�y+*c�Ak
��j�7p�,p���`�8|T�0����A<0BG	;әO�i���`�ѯ���s�{z�u|8���V�&�&�=s�A�k�y��2z7�r��!t��3q,��t�!�Dz2(Da��JH+F�Y�r�V8�����c	�n-MѸ�;�s�`1_ck���dwi�a?�����u�g�����pr�ʋ�y��,i��({ 㧂��sT�>��hz+�r�7�@�����iU�E��@�R��߽�$%��A�u�66�g���%����2�g��a�-�<��k5Y ��v�Qq2ύt����{=�1u�K3���RKk@�-Y�r�^��$$6zJ4��G�@�ݨÈS��C\�Z�nZ�,JT�䟪q��&.�L�S����d��Q�����$���,��dQ��9Ԫ��r;\�E�o����'��Ee��Ј�u��|U�~!�����+N�| ��C~bǞ� �>��򭅭ӽ6*K��|f����2�m�g�"�:cZ��4CRZ��md��u�Ӷށxo�x5�����#]k��~���)G�N��9�q_!
%Y�����V.�u#1��*p�����k?�h�:�Mdؘa�Y����Buy9��Al��m�������|����͔G����e����Iʟy�x�x���}c�?���z�|��=����J�Q��)&"ڷi�l��<
 �iu�}�Ixa��5�E���(I)H�'N�yR�L8���|DC��_,.����&e�+1˄{���#�R -���A�j8�8 :�Y[�pG���.��2�\�6K�n�m?��p�Y��?Y}Ӊ��;��}�&�	��� �n�!W���ֿ�P�-fO��q�u]��"ɆQ�@ߴ�Q��2�$��'1-�O$����9�`�r�-_Q�s��߮�̳����(�Tؾ1P��<cpL�~�q�X�sXfQ*�1.���e�i�Z�>#�D�l6Ub�<��W �BP�����5��EH~�Hf��n�ˉE	�6��S�7<���G�*�Z��@�GgI�Iw(�a��$���]JYsm3���ZFF8�3ɯ:O��v����ܓ!�tA��e�K���<:�x%9}��-S�SΕ�,(���%��`���k�����iCz0��H(�IH�2�zZu^Q}�L��RM{b��h���5�-�0u�d��P�<`�������g����C	v�����繾Gual|����_�6������K�>����(Aj]�5�R[z�bf�LP\�:�ϣ��.��TF{�^��x�Ԛ���4i���v��+���n{+�᝘�S����<�rD�r1�}R�JpN�){A��hb\n���aD\�B��y,��ء���|�H�gd�_��~�_��^y�mXy}�	6Г�
�.���G�U3�H{�H�FT"��^�8�,��}�&ϭKsx8e�"4[;��Z�QX�>�n��]w!��w��D�?c����<�n�۬P����N��p�Q0,��N�����q�~6�_�b6����e4��k����RP��[�n��%��#��^oB$��Wب���YSz�lE��ۧa���v8��� e1����$��%q�
��ԥi�?��C~ĩ��Ti
Ut"�Ӣ$��Ǟ�:�^8P���.�uz���E�\���#��a�!����b���cE�!���K���Q�d��+�6*0O!!�S�9E��LW�(�3�8�Ŕ��BҸ��+���2��0!��׈%�~��5��
�o��2��wް�J���(�Izd2 ��.�ىP:b�/vj�p��ɓ��_���%S��+�u�S�0y�E��i��#{K8�m�M^�������x�T�?���J�O�N��u���c;Ȼ�W^�I^K�u���p(g���%��*�U=^�}���^ѣ�+�I~&�LB��ʎ�@�c~7�����>ه��g��H�`A< ��t�~�2�������bY��c^v��͇�t�x���3T,2s (%N�7�E�Fl6�t��E׍[�9;������|��������!L�ơ��� 4	��R1d�H,+���c�Ϡ����ٯ�hFr�B�Q2�v�8�!^b��m���f}Mj�Q���da�$ŭ�ɍ�*|�KO ��卺a�P���t���+��21�y���E��b�:��Ep�v)��/��1 ��[[@T4�N����J��}]��L=w�D��o�>�Z'��K������9݄��]��5��>����y��1ш�n�z���Ӱ{���RX���ý��n����X3���F��k�5*U9ڭ�9�큠��]X�9�Z�֓�s&qQ���J����6���]!/�G��@ux(S���Ԯ�q���7z��s
�vC$6kT&I��F7��'�ш���{oܐ&2'ȶ��10U������)�#I�>�.0��kd�M�x� @r<�N��Z-9xw���g�����dØ��(*�7b ��>���z�3E!��7}�"��b�fkֱGW_4V=��kv.�T�\�֥0k/��H�`�[[ꩿ.8���$�(�m�zg>�/{���HM�&f{��#+���!���(�v-Ѳ�;��&�5ft����<<9[����kfp�ke��U�tɁ[�6-L��<+��=^gIB(i���9Ψ��/j؉�4����_�b漨�ؓ�w>�֫�;[& e�Bu:��E
�\��u���a� �g�ls��T�)1�&G��'n���9e2��3w?j����a*I�wuh���-L�e��w�����P���'G�N<�	�����Wb_B=k$kG��gPY���_S|��Zs�J+h:���Uռ��3)��N��l���&ظWOh��o�ԧ6�1ʙ�o��y�_�Ұ
�V��?.��Ҫ�Nf��Z4~�b }�0��S~�t�_)i��Ft��V��5$#���Zl�
$����$�TM����zy0�������T�6"ۯ����
4MK��%���t�n,w)�w��f��㇘*Ķ�>�E��uo|�"�p�4E���=�c��E��_vlkOʨ��m	��պ���3U�W������'|��9�~�FEU���s:�������9���uX�/d}���������쯩(P��?�H����Aqf��McV��n�*��y�%�SGe%2,|`nOc����G���=�q�aZ��Ep�!��x��i���� 8�]>i���݋Ͱ��=�j��B��4��&��b���	s}8G��V_�s,��������hp-�����GyY�m����5��8���As1:�1�i�V��G���2�$�;֐�����}��^6�t���z�'G ǥ�����E�����?���*���n����Ê�%���s����Q��!�!��3�Ws^a�@J�� A:U_Ɠ8a@�x[Ѯmi�F-}ef��T�{�t��/.$����)����aZ�&n�H�� �LP9���W$�8�d
����a7�.�Ig��yC?cJ���Iu"�.*2��|X弴=�!�:_����>��`?M��z�nHq#+{ ���h����gB��Z�����T�'��0���B��߫�X��[�%M,<��Å�8Z5lپR���Ȩ������@#{f(���J�5�&�4�>��.&֍\��E�Ǖm���1VT9Bc���T/>�)�&��T]n���;�S�iE;�,�@5����?�.���A�ҙ�u�ʆ�#����W�;��+kQ1��:�~�6����\��^�)LNc>�m�tl�Ia����7�}�E����,�� TOG�X44�k~G����������C��i���U<{��z7�;�	'=2��q]�>v�|ωXz� �Kz��!���٤ifC�,ɰ��2�������iB�& F�O`� ,b�݌R,)�Ǩyu�;�Gi��՟`��N͠����
�*$GB�2J�Iԉ ���+)�:+לQ�֦y���F叄9�Vʂ��D�vb﯍��P i�����X����O?���Ph諘b[�G�:�QU���+�ɗߨ��4�I�t����.j:����\gL]f���iYd,T0�4��2˧!�ڵo�ʂ�*^3K^�e�VB,���[Obkon���Y�@�^�����v���fW��5���ߖ%�;`Nr��4�D t�it2����J���q-@��I��G3[��0K�+E7����3HBO��{���&r�J��dvc�06`[u�ɗ�d�F�'��.5���Q��