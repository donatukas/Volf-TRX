
module DEBUG (
	probe);	

	input	[23:0]	probe;
endmodule
