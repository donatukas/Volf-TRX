
module DEBUG2 (
	probe);	

	input	[2:0]	probe;
endmodule
