��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5��¼��&G��ˬ�|���Z���7���U���xo��(��g�n���p,b`�fC���ǌ�n�g�m�t���6+��ݟ���Ki�e�$��.�x�/�AGJ�����`��E7��,����Y@�:F��� = ��3�����9�i����U�#�i�A�)}�,|7�V��&��*�IC[-'��Q�.�۳��"iy��▇53}أ']��"�������ۅ���[��gѷ,�Ash�_�kp�5	�ֆ��)�>U'q�7�s��搖�u����6������P���߯����o|�Kl<��E�F����V�l�Y�ET� �y�&U�c�-�j�4%V=�][������n��,}ݞ/�*w�2hz/��'&Ì��E;U�0V��'uq�"Uo�ғ�d�BH��õ�a��}07I͑�
۰�E��*��h�'�@Й����b?�T�����b��W�u1k���˓�;�/���3� �K���Э82����Z"2��>�������Xn���Q͒A���v��nPS;=�\{>�t &l+R3�#���t �J!��AgbC�T���^�-��^�����Y���w���=yp9����t��vQ��J;�=KH�k����,JT���������a7Q.��Tc�O�zB���_G%����>W�6d8�cZQc��
سϹ���w�����ri�OB�t�?�m�/|��+�j�-��P�G�'���TxQ��P$��40_��UA)�x�3�G�6��������%�C��^x]߆�~e���d��k����i�}��nƏ5{��. L�Zԓ^�����n�oJ��"L9:���c����������H�D�)�n�	X�Ux�u� ?� ;\��Z�\���t�?O�T.�90UR%I/Z��������v'�+ࡥ.�6�@_�=���
����n��+�Հ�?����+@������kE������<��ɹ��e���H���OM����úJN2��A�
���-��>�yu��F�����wխ9	�8�UUǉ�I�vFʐ%7�A���~v��������t��Ls���)Օ����O���2�{�Ya/��{�se���]ƚ��ܵs�@˓C��n'�&��j1=��>S�9C4�	��*)P^f)̔�"����}y��`}!97�wa���QS�.2�a� #�V��U��5/a��|��V�� MA��;E�B͎����m��O˖-a�G�a�Ӱ���]��*�A?rv+��Wk����<�����s��Q0��7h28�f扛~�QM��8����^}�a�����Sq��ڰ�f}�<�*������C�|�����!�d�����#��M#�R�{�V�[��J���R�`�8qY��>����`��L	�w����&�mBrzt�(�
�/@t V9�U��K�x2b�H|�C�p�D��V��i/yU�Q�͐��@a7�#t��OX�0�����(���c��3��1q��Idn��։b�U�Q��|��N-�\i����\�s�9K�7|�L4|��s�5;�:�����ؖ��RJ
Ƥ�|(��S����i��$�d��	G�&:���ϋcz��oJv�����NL��9��b v�10�6���Rn��\b�mp��{�]�Ȥα�ez�;�9��Q5�e|v�fn&�Z��-f�+���o�_*���k�N"c;}�J��9��q۩%�c�����@r���
gDN�L�r��%�c�hD��C��<}�,(��\��R��;��["+�$&�N�n�伯����X��
���X���T�.��-�;���U��P�J7�k]׋���"�am�L/�Q�=n�S!��hՉ��Uo�j� � ��2P&���U��M%],�nn
�9�5Bc��5�|�&θE��"��g����\8�W!D��S����Ju�D�ȷ���z/.~T<k��o���3}����%]p�٭Yo<y<������]�(�����AU
�%�����Uw�������K�/��`i���gQ]�������K���fK?���o����`��@�$�n!1q����}ec�a'����R4�H�:���n};�H��,'[K��Pg�G�3D8҆�Q>�~�ڥa;3���<����l� 1ַ�_	-��t��˖@��3`�0��H���[�ik�̗�a,ď.���d�)�y�ld��?_������Eq�/���%<V�>�]Yi������*! ���	���3T_	Y�<��3��\@~8�5따��?tR�<uL N���a�g��2��Oya����U��|�%.*�6/�Ic�����:�Ab����L�|�F\��ʎ��8Y�2]tP�W?�BL��1��G{�*��E۹�(���2���*��E\4�a���O�	�{�=Z���
�.�0����̴&�gGe�z������'���޷m�M�X�<��En~Kc�����v�V�ZQejj���=I����rd)d��4�K�h�	���+�FJ|���E%���q6������
9:�E�?-Dл�A{1�ia\!b;�,�1w�2|J�U���v��~,����[J�cq=
�;�*P��*~URG��@��G;�e�G�s�v��8�6�@o���QS�����������v��M�[�HuF�n���GӅ�}���YH:�Z�%Z��?z5�w�f�f���(�FS���#BC�/ ���(�H���#�;��|<�<��=�䞳���:�Y����[	����ɉ�x��Ĥ�5c���8��ok��h��6�O�৲b��Q����'�XOA�v�Lu��ű	++nGΖ;�3�RY,�B=* J,��&�A�DϫEi���aAYT�#��)��3��?�A_#U)ت��Ь�Hկ��2K�Ѭ��"$��1[9#�*`�X�d�C�C{��#Nqu�0zШb�搬̩��U�[>(Y��?���f��[K޲N������reB�a�J/����%���q�c�I��K������5�i{9��{��F ��ƿ��s�S�&�S�D����<��X0��t��1��2�=Ղ/W	�:�&��`v����nF��U�;�=���:JE#�]�uS���<�5^N�l:V�~h&F+�KE��Q��n�-r�T�rr�N�Dj�f`g6����UM/*4Ճ�'�sannr��m=�g?Y3r�j�L��
Zw㭨���8���$C�4Ap\H��Î��hK�۽�G�I���1����6���J�{�V���\(�C"u5<�*�Z�3f}d@Z��b1���!H��ԓZ�b���(����i=z ӥ;��7��4���m��2JD_04z\��zhixII�.֦�[������e�׎���~��[������1?����/��qJ �!�\X���X�S+�wr"|���IQqҨ�7�f�QVs�������0K���?�zķ����pߚ��8����!Ư/5H�A�%<7�|�Xu{m���'�����=O������ KH�	̼��g�v��ezSx�D��$�(�%�'-7.A`Ͼ�׮n]>����5]t��z��nw�O&���b��Ib'J��9)R� ��b�e�V���ɨ6� fP	�إ�c�0ǂL<0驇����"���0�8�}"��U�3:��Q���63k��������l��\�҇���F�!0�	��2q��`c��H����1� ?��������税��9C�7}�}=�턯³02�*�q�\�����)�C���5�>�jQQ�Ad/Y.w�I��?�V]"�j`�dK'9���� ,ғ!:�Ԃ� ������Լ5b�WP�7<د�5R��ъW�}u ����qؓ�"j^Z�	g$0�F��j,!�M�ʱ�����aH�gs'�B�K�U;�ҏ��k;�U6�[�,��?!k�RZ�
�a��¯���E��v�)E�"�Kt�^����v�}�0/4IܿQIc��`:��7D]&�cu�^ݺ�:&6�x�o�d>UAi��Q�Ʃ�S<ZCd��S��H��Su�I��F�'M>&���_���:�y����#��N���%EB�`�^��_�D�[C��C���G�^3�)��s�!�_E"��jN�����aRV¯G�?&���g>����a94v��-�>М��(���UX�d�\B���o:�s�