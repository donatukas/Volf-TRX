��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U<-T�M��e|6���0�-���Zu���ϊ���Q�|:g!�����`~d��ЖU��BJ��U���)�   ��Ħ��9�:mF6!�E���~`0��I
�<�?hHOW%��)�@5�N;f�b�\�'xyG@��ҭ���*ʌ��L'���&����n�x��+��ę�߱�g3���"������u.�6Z���vٸ��ST� kBE�J跄�'GDXD-���hp�UBʅA2��??�1�#Q���/yG��;V*$�e�'�ǽoZċ38��1��5��{�z�u���H,Ftd��6��b�����W����� �3��/�8ҧ��A@��3[d�0:��+��3=�$�Vs�8�(�t�\���z]� N|yJK�~��+D^yu��>�!�h6FِVD)	q?�[�������6-�؄�;C7�,�
��é/@4ָ`�uՑ^��u�IÞ��U�}�{��]@+b����B�(�{�bF�U�fQ��l�L�̀-*6�}Nےоo[z���IC�G�.���\0䳂]@͗�E�~��|��be*����(렠��Pd-yg-���ԯT�ċ��N~F���S�[U���{��ӿ��oaN0"�q��ֳ�b�S @٥r�ir�0�'QA�!�M�\���Q7�2?@�z�y�]��s�)B
b�^`n��6���˂xD����p�5�"�l����d�� ����(���T�3O�6$u���{C���E\b����j<>�4�Y��za�n�1>3��*6��.��[wpF��#*�>�}�T�C�������#5{31�xD��=�`������d�O̒M��<�'�b��3g��׉��/;��Q^����0N7�N�5��Ҫ�g�̻���K��u;� �d�uI�>�|'l��ČͿ1��pdo|�V��r��p^��9^�f��͹�B2ߛ�`��~�����w}�é(n�����߭@9J�mgǀ�Y1�F�`ө���Uڒ<Q>��bz^-%^��r�ߠ��>fRXr�4{]�j����p~H��]s�/ �|'&?XE�n�c��)
��t��Fg�t&�A3�+������+\��+V�کP$�FfC��5���N��ʝ�+��c�Ԃ��%��Y�?j���đ���2"�W�H���CUd��m��j�b	+̀�ӶpJi�!�rl盼?B=�1�\ҽD@O��'6�tИ�䟼������GC���:�E�W^q�|Io���D��
&^�./	��M'1[�Z �"і1-�UŤi1	ۤl�~���}����A�4]���M��j����
́ȟM,E%44�w�	���#�>DX{������kt�di�.l�QtSi_���b^��b%(�2�����[��#뇙����I�� Z�-�/s���bu=B�	�y�_Ϭ0����z�*}�SOb�k+9-�xp.�TE�~-*;3�}຀��pŧ{���	�h*GZT��(i�Gb$�X�I�x��8?��p �dt脇�2��t�|�(�4��@�Yb�
�)g�T5�������v	�o��
�eTA{��XӸ]�'�.'��#���q��%>�=�eہ����_�����<j����u{�P���])�\(
��aj ʰ|jvL;q.���{I\�$;�Z�z������K��E�����u��tf�nC�أ�6��هZ�J6�e!qO(Dk���ر����G�o�]���>8�4R���S�Zrl�m�G�����R���6Ɩ�-�Q��J(�p�q�x<��l<yo<`\l7
pw�����ņw�̄��pab��z�dy�R�2{�@〜��DX�LV(]�s������ �w��L�]�;�)4�e��`�A<5�g�x��gNc��*	�q���.ر�!H�Dg!���M[o�p4&��~G�6�����sM�	���-���<��i|���B�K�),Yu�i&�`�z�8�>7)$4�[�����&T�u�S6��ĉS�F�U$"	�h��`��gU�(�Tj����ܒ�S��o��{�0�F�g�ܐ�ˎ�L@J�Rw��"�075����Prt1n�����%�O� �G�J\'�_;#H�l�����t��I�w��}	�dAA��z3Q���X���2ɹ}��XN$3�E/�x�ۊ]�Σ3f�q_�S����x����=�r�BU�"��7�;ػ��`&�i��j�<�a��2�����jh� �$&�[W�Y�XP=@>���O�$��eÌ�Ə7������'���}v��V�|x���X�UC��4��������t/���8wD�F�:��k/B��Wۑ�������D�1Ͱ�@Q�u��Z���*)�X����&e	�����f����G�	c�&���j��z!�0�� ������O"Sk�C枦�\��m�0�ӣ	����4�<@�h�Fq�Ki�瀧U��^[i���f���}��<M�C�q�F�
ͳ��&@(\BKejC'�L�g^,��.͌tfI�I?O�	0�E��W	|�s��n�ƒzz^���Arp=y�C��=�Ul��x#�V`]]�8Gs?���ԙ��C��]!Y���0�N�&Њ��_+_R*�t..5tL�OgX�yx�nǪ|(t��ͯk��?\᚜��x_uoBb��K���gJ5{@�)˩�x�X�IvC+Z�bE�YL�s{��8����:n�x��uf��:��A�b�����n~���j��bm�v�f��,^ϐE���|�EER�?��B��.�>�����, PZ�|f�ՙ-�z����~^���.�>��Đj�b��� �`y:e�H��Z"?�x�����4*��@��_�~��T�#�/��u���o�����5<AP���
�q`�/�3x(��+�##w���h��MV-ݿ��E΅�ޖIÊE؊�	���� r�Q߈X�.x&�uJ%���5�tt
 ��9{�Pߒ��������4�z�?d���slDe��EͶ���~��ڎ\��Y$#�yl�Pt:t������|݉���,;������ܶP����ut��Ö-��Ϳk��"	�L��[;-e	���Ԗ1�*���������SkV��m8h�&�&1�|D��VI턽�q�r�Ov���^ji�j�����y�h�׷�ᑉɅr
��d2Q\>���*�-EH�{G���	49�i�Ⱥ���%I���os�:�\�j��wA1�E��%&�۰wf��P;<��K���^`e���g��D�z���lol�_Y�i�h��E1�yY3���2˻�va{n��d�x�v���.V�9U�3��G�}�)�Y��f�MΆ�E�,x{�v�#mH.�	zbc�o�����?Q��ל/ �������j#5�c�#�v���C�課��I��V[�-�՗��林�ttS�,��L��ӌ?AH��~��b�D����*��CB� n��2o�*��ˡ�J�L�q!��}5�I�r8�80�`32	�4	8��Pn
�].S+����j�o��!G�5�*1VX*�\I�G�"�s����Q&�������!�j�pV��$'�@H[vx��\o�
��� |S���%�?6���I;�s'��4�����Hd�;�4�H����/J���d��s�����f����p�p�h�����y�ړ�#)R���wSLf�6E
�7W�i�M��N��=�C.���Dφؓsa��o���Q�y��B��K�6��}�����)W�;+ʒ��A�-��@,zyU�Vm��	Ɲ_��o�,)d.�����P���W[{���� ����k�Ũ��v�((����`XŨ��O�e1ܟW��k���q{U�cu��.���0k%�2�xQ�:k�[?V[�g�e��_�o2P�(88���S�������-���{kO�q.�$�r�9n�@���!�c	.@����t
�V�rկ�<�YV�����C���r��^���ʵ�˶����2��hn:�zN��A���Ѡ�1+5�8-|���R�j���y{,���5B@���h�<�\�H���*w2s '� n���(J�k�����橒+��UiO����_�J���41�we�-3��+��`���ܛU��(wx-B8��X��;��/E������s�oK�&+{Mz��$3��^#u���ڪ�#�cƽ��9��˶��5
_`A$��#@��y �����1"N,��Y +q$'4�"?��)ȏT�����Ye�t�-Ϙ~-��u,r��&��TrG�e�B8g��
�%�$��&j6���P�F�Tﭡs8=�;�M���o�5B��������f�Q����N�@c���)bj���"H� �0Uj��X���]�8[z+9��,��p^N���6 e������-*�%��]9B�m�ZV��?��]��V�9a�W7���#�DҭrG~Rd8�1���'�@ykP��������2��`:\��3�O=�8P�-w8�ET�G��z��fAr�-tʄ˦mq�M�
��J�Htb���槹�:���y���$V����CD �ڞ�>�k��8X��M���3��ڠ�����y�?��7�Dm�v�����b-�ۗ�;��CO�]��j|�g��( /�L$���iJQ����}�֧��	�/��^���c�]s��~Ar��Lt�I��T5���I9O(t���<��l�L1��F�*�ha�sE �c�\�ז\4: Q^hf�� ����ȸB���F`���<Ons��<�K�9Z2�'a����Tw�t�
�?�ƞv�>�#x���<
[��-����I��q����-��E�b����yJ����r����¥��af�!�OAQ�OS
�-Fy�%�VP��<A"�[�T�9���~�b��[���Y]}��Wn��8H�AA�ɱ[��7M�ywh<g"����p�.
 z��,28p�"71�Z�1o_Tj��Asu4�j��16��u�J�_F��D;n �g��Ƒ�Iy�i��@���vi�5���Wn�@dxIJ�$��~�4<�mr���)rym?A��17��z�o��3��k��j��nM�i�g��I�ȹ�0�_�F�T�ӦsY~w�^�?�� ���z����"�3	�?W1�D.N�#��a_��'����,MoAWg)�����k1]6AY����rab�x�G ��H�k :�t-��]}'��ѳ;�(��:�/*�4P��� �����|�[9�8�E埣
07Y�e���Xe� "�!�,<%j%jUC��}��Kvz@������;Ja@����A��@稉�ܲ�E�>���jL���I���'��=3B�e{���7���*2�qwY�=�T�uR \��Km��l�Y��f�� ���Ձwli_4O�5�����O/���	M�p��gQ�s�p���Ϲk�qȵ��3qDM
%�����)�9��g����]v���!�����[<\��װ��>8g����g�:���z9r~0�0�T{,�G�(�MD�R�t�_�/�m]��ѹ��S�r[�KM������J����R��FXva-<Ff(�.�gj��e��lt	��)4��|��&RFFƻ�~ϯ�F��L�ɜ瓲oԻ+�` �/����6�^����];C����n�x�y�aԋ�
a�Q�Z��6o�ZvG�X�N<��9@�,��ǦF �x�ٗ#��}��~���݊�#�1+v�S
��3%����#I��#����q�&��~���NmjCѬt��#P�llR/���mc�$VmK"�e��3n�p_��Rb���u�[��<�$Q:�'h��;Ǒ�N�pJxK&T-xË�F*��d�C��
qZf���j��_]�y�Fjlٷ/�����6t�)~�c�wd�;1��k��-�*����� Ҍ��z�"�p'ڌ������W��q�K�|(�u��䳮+��p�8aKX����q<F;�u���p"$|��h�D~
Щ������HC�c@Z��{���'�^Y���D�f=����5����m~�#���G!�
Ĭ�j@�`a�m��ku�% "��po�2��d�"J:��&�����M��п�y\;���WE՗��8x_��_�{���ƉǬ��fb����[DY瀻t��0#������-�. �V����R�K��уp��]�};ߚ�R	��X���BS�ZL�����Q����S�Ȼ��zhu�U��E-���z,5�WK�� �y~�d�I��J��z�ӯ��I�*ij���ie����B�[)�E�)�e��R�|���^o��&�����	��;ԕ��(��r65���R=��B���