��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.yu�=�6��MYN9dI$s��z�������d:2�p����?4��==��*˜�"}�h������<V��� �넨+���)ÒG���(���\y��$����@��J���Ք���|��~� ��͇y��W��^�+�r���<w�T�^��}|K�����?������w�He��<g���8�9{��-Խfa�L�
�@����U���q�2�.��W�禝`s5��$�.(�Ҍ8�Í�y�y]�0jx"�6V6�3��fe h!��()[yDsr�(IF�r�#��#Z�.d��3��}>������-e�4�p5�VQ����-�<G����f�S�\He~����E�)�-��0�"]�P����:��~����]�҇B�=�m���\(N����i��Ӱ�v��Q�Da6�1��5ENq|q�� �����*��x󄬉�.�^��~��,@�iۍ&���*�~3F��[nE�.����f����~��Bส9_֧��/��f�j@�F�]���Y�D6���l�R$���.�;R(���&ّ�����<��j5hf�A���H x�Y6�m���z߬k3�T�)/ܠ��a��*�ՏhN�P |L����40p�W*�l��#�Xg�]ݔ�<��" L�.����$+�B���^f�)�Ғ��'M�p�4Q�+3�y�r��XȻz���C��i�w��v>bڠ����s)���a�(��3����x��Y��h�]tn�,��.���ӄ�GSl� ����˓������k��_�E9:��~��:��ʻ}��S�����oC��TŢ�ʡQ�%o���_�2�BW���u���{��^v��-2%�c���ߑ�P�:s���Yհ$sVS� �ʝ6��J�YB��H<Y���M����b3��F��Z�A�>wv��:������lgk$ΜI8�I�%P�QH~�A<%��_W}�S4�<P�7G�lJߋNz��r9i�W�*`7���K2SJ���V�z���Tm�n{�gXZ��M���X�w,[M+O��j�9q˹2��:��i�'�%q�ol��@���&��P��d���
8����	���.'v���".!���!"�݇i\ʄM��
��f���RM�ad4�4q�����NǱ�"䂃qpU����D?���DBt�-�yf�N�;�C��W�\�Pz5����j���h�5 ˴=[���R�����<���S��mx�*��
��?O��;v�̶-�Ʊ|���^����v���l�(g]uȣ�;uµQ�yY����+?H��,�r��� 4a�I��k���o6i�evuv�4ﴝ���K�2�D{c9H|����[o��Ђ��B+&}����D_��)���"�Zn#��L!�����#�Ɂ@ S��lT���]H%���¥�F�!��4�(9Z�:C8�
�J�^w�b��^�+������H��=�^�n#��L\�헹o���nwA,p+�	
+/��~|�\��j���͗@?���]�����
��&�t���=)������N���b	����y��Pq���a+3#Z�󚗑�k�H�a"f�(��JA��
�Z� �ؾ#��_me�ʹӽfM�"0���YDQ�4a;4�2ʥȸ�ull%���탻�h������0���3�#������DRZ͎��A��_�e萕���J~��HA�L��A��'����

�*6�@њ���T��e�d��f��ŘE�\�۸��k$�:G:a�(���8��ͻ�~�h���G�\g��6�n���4�jQ�X��A��"�&�G+�x����堌�p9�x�u���T���L_G��)��7�D~�X�Li\�ᯯ]�iy�Ь�n}�,=�������N�n��N&.&�ĶE���@eK�9ҫa;�&�L��zjZ�敢?�����X����"��O���`j>�9�0U�%g�Ch:�����p,_���ٹ�VU��@�b����U�)�-P��L�[��B�����lѫ	��+
f ��RЀ8f�d�:�4��[���z�6'#��d�9G
R��U����z�`�4��g�w�<	��͹D^�ݗd%JMN%�#������Ƴ�:��S�6ڰ	�N(c�%�#x��M� \��9�M��1=Q���Y����ve�%a����𞸃Zt��NfR��49��og�1怍�}�od���$�;��Ӎ�Hb4v_"�>~�lu�s$ڿ���l=��) �B�|�I�!���;G���J���<�[�'����~�e�Aj��\��)k�����x������|�GX2��fA\x�����C�}��i]ϳJ�S�Qgd�Y����r�N��$��
{�t^U�cm�@�^���`�,KEf��mb���3�i�1��a��9�h��]���'7�~��Vt��ܒ�M ُ��/z��Q��Cp߿�}1��5~e�l�8R�2&�K�AȾ"rbf�T�f%��^���@$��
}1h�5S���0;��NՔB�'6�㣭�H�{ls���(���o�Gb�X�&-�(�vN;�$A7�ܞ�ns�w�'`(dlHaJWe��k���ʌ�ȯb"���- k���������B��p�������6��b\����a�V#	�7�;�X�\i(�Ɂ� 2i;�p�\�E�ɌS?'fst,\�/� h�G#�F�V���"�5)�GL��y(5R���� �!� w;�`�	ms݁|u/�/��9�*�����ӎ�XT��{Z�u���c��aW��Hѓ�#[�m	g4|�r?�S���ǀx�{�mMt�^���RT	<��_)H�^����jrż	���KwȉU�ܐ����g�s4c
��Ň]���@E�������f�_�G<mG��j�RP��.fڬ���~��[2Jn�?!��J�U�K��+I*��	ws����j�-բ I��e�Z��lإl�࿆5�$`[ �O�	vɛQ������`@M�D.�9�{Q�7��͞蔯�0�9�85y�v�OEU��M�Cl�82�l����zء�A����J�_��o��x�����Ǐ�M��R_�짣n�lH��VV����\B���1��\�L'���!�ƤV���]����}�]�PR=�W2!�r���5ZwXh`}1�%4Xlm��1�:�
��O�_��A�ټU�4���/�]�1% *q #`�̣�b�/����nU������+=�Z^S�^J΂$�\p�B�Np\'ì��m��P��7��u�[����o�f�7,cf�zٗ�D4�c!�7B�?��A�6�#��(�7���ֹ�g�Ȥ����h\����P	vZ�o�t<� �������,� e�#�+Is��u�m�\n˳��1���<����Ƶ�KH���q>e)�=z�ڶ�A"�Y���;C\����U	[�4�'2�U��22a�z�]_;V3�-�&Hv�����+n=�O��)�+���@x(	�w�i�����}�B�=�@i��P�lGfj>l��sT�ڼ<ed�g
���B3יi޵��tB�5mI(&GA����8l}'*����M����_��q��!2V�S�1p��l��Q�(��K��F�8]d7Ob0*�ݐ���q�B�_JЗG�=ѣ��(oZn�sv�a%�R.<�#�\A���[}�OV\��߸�r}�߮�C��9 T2�..@�5\��b��ц}��IT8�uk�Sp��a�=ׅ�HWz���hN�H�H�$��-�*�?�󜦥�ʰU��{-���)���|U����-���$�_��;O���x�U?��#��i̇m��IV+P�G�#ŏ���o�pNyӗ��r��k ��.?x�KI�$ef�u��� �/���ӽ<m�G���0����g+�� �Df1��o�J�'n��%kk�sZ�گF�~,bB kM·|���C8�ꙡ�eu}A0b���Nij���W���7��kд��;�Ѧ���O.D�̯������aY�w�]`��n���RL�����FR�tr�=��Ί�(�?C���f�`�$���G�����I���΂�x=�}p��;�|6ۣn�	�c���ڸXF4�`����Q� �p~�8t�:�c��jA�7�Z������4g��xF`]���<�#�p�@Q#�:�b�;�XB>��z}B+�RE]|95�`2�7\�璵�#2q$�
ԯ�E,�S�͍��dN�?�LU0fLܪiڨFcv�Z	3��֣��?-��o��"��U�'���I�u�W1?�h�W�v���a,zx2qZĕ%C6|�I�DG(Pޘg��T}�:��p��� ����Az����r�B�5��Z:I�`�R���Jg�{{��,��i<z�dɛ�_��>�4m?Gӛ�'�¿�����&��N=�zM㰜�ů����3q;	��(#���E&@�x�E�0!�%D.#ya�}���z �4i�dA�����OX���%�~�[NH�Yv�Kt�z�A���X!X
��TفM�:ש�MH��)����9��s��u��)Z�r���[��r�$V"��m�%.[��{��]e�����m�x�*��JK�1 (�3�R�!i��R��A�"Q�v�gK��'S d	H}6]R ���&X�z�ӽs�-l�՟.��g���^0�qDMo ���=���y���-0�p������#c���Sø+L�lhIҞ�g�ul�KX�I�@�~�V+���L�Q�"7���f��ˣ���ه]8�'����y����7���^�(7*�To�8�<��ꏵW_�D�-nE=l?�����q�����9�12��y��R	d�ʊ�+�3{.�mr��5q<EP�0�Mo��q�a��i��}:-�]AQ$���ݵx����S3^���6j*e��B�i+i �<"��\�;5��űa�A�gc�/��'5_VH�����n=�;�?2�]
o�^��%����w�������x0�p�@�U��ߘ��Rg�����a�|��G4�ˁ&W���R��y">o1�D���J��S���C�/qSna���d�,ϖ�c:JG�h�m:�����Q���c-\p|��n������3�N���X\L��Ml���P���v'�k�"����)u�#㚶A�M�W$�<"��恕�\�4���dR�3�y6���B��4��9:;�MV55.���?r�1�����sq��3��Z2��`��}'�iUj~#���	��}R	����BI#�%�o$�@&e����W�Ɋ�QB���m��\-�̣��1�e���5v`�.D�8�����l�̿ƅ�ke���t�H(��)�>�\�+�8�Ssd	���Wx'�09���>���Ft���V�,�g��V��d
�Vf@tŝ
akƽ�F�ɯ�(Yn#�����~PϜ7	v�@���W�,���j��bR��ƽ�Ua�E��m������:u(�42��P�e�ۦ=e褈x?���z��9Ղ����)��;
��_�#zFYL�>w&$ӚtS#�R��]������_vQ$ZE jώ������w���6�,��z������n|��Oy�)�엵�r��m��Y� r+i��)<)�%�#����}5 �8w�%��,#�F����;P�{v���2��������� �l��Ԭ��'�?��C�<ޱ�v�K$.��ՁNj���f� �*Tl�T��T�C�N�Z�((�D�%��,=��J-� �9yQ��c���^iG��,�
;آ!�<�.�d�@hҷz�����ά�� Xkx�D̎�$eX��1�o�ٺ���i����{A���Be1ي�R���j��42�����Kyl��KB&g�>U��T|� �F�wA�n�yN����Z��	�����������0;����@Pg�Z.]�o�A�,�9��b����G�$�%~Mj�>��Q�ܹ�;�K�
�0v_)�Z��Z]�Ɨ:�ViCn�::�u��9)DO
���!��f��ǔ�a���ǌ~H$�z#x䵩���_<\��6�BA��"�3��u`�����"��KfB�4 �¶��Uc��11Ci�+U���󼠹���)�����2�/��g�?A�z �ZZr�>��)E:B7Nk|0#���j��ޥ��������l�š������d_��������ST͓�kS�%N��!墦~��k!�o�����!F"��{�t��>���
t�[~�=�v�e�d��CІ{9gw9�s{��$�Os7���Z�/T��uu��~ɇUD��{��fb;��C��k?{<�ec ��	r��h{Kf��x�)~��w�E���h��CL�'MI1�P zn�{AM�����-���|l���*����>|����Dk�<)@K�r���FOضX�T��Ӿ̶��J�BzOws�V�_����X�4�
���tҽU(����b�����3Xxҥ�g_V�*���}[�Ҁ�v�L��<YoS�8���Q�,���rs|B6�Gv���S ͠)g	_�T�����F��^�}�}���DZ3L;41NA��i��̲�b��u�}Ϻ�p_ى��{Ļx��D��-pR��H�<�}UxL��C��s;�/�\����o��4,zo�`����2�d¯�ծq�t��Ӓ��``8�.���Aelm�H�N�'!�j�}0�-��"n�iC�<ͦ7p]���i�O���s��vSj�D�)=�|�s����tqb�/�\W/`
V��IP�[�xsB�2�0�8>31[q�{_�
b��bJ��F���¼����m��\�APn�\(3+�TۖiXRsX�̑�p����s�?ɠZ|ͅ�S�m켒��r:�:�C�K�����h/���e<�f���96ߙ�b�#x�ػ��؛?;ˇRyZu�\N�~��r����zg'u�y�M#D�&/�7d��3ЬoJ#3�3~Bb�0��HG<��%�x{�#\JLMj�c��z��6�'1�y��:T"/Dg�0Sx�Z�҄�k���߶-��JDuu�j�w�"D�=F�����V��&ɫ���-��P��ن���}��.<�w��u�����;s�_!��J������0�(8V";pKt�ٕࢻI+�6\&����ج��kX6J�:�MD0���qsZDmy��0i�e�R	m$��eg��2�fl </>��5v/{���?������9҈#�PXg鈞��X��:]�o=ǝ�|��
D�w������+�L����uL�ђ��oG��X�w�޼�Լ��).x��o��gN�Ƃ���׏{�!�c�>�-]����,cn!YF�>g`��̈́w�w0�Zmqo�����r;��F^�+�����ڛ!M�u�	�o�M�S�����'ʇ?��J�s�~��y
Äo|x�º�	J�Ә6��rt0JUd��T�1����
��������7��`�?t� �%X����M
r�ti%�|	��A�ͥ9�u:�
5���Qiɏ�a~Q�>�]�G�D��p���n��9�Z�����v�� �b��J����w��-��C�#8,x5����"����w1<G+E1J=Y���M�;��MG�0
��AfǮ8t[ �b�N�(�/ �RS��Y#ud�9qB�F� ڍ#��Bjެv�ܲqu0P�+h��O��[��&j1�}�ֹѐ�^{���p�Я�D�~7���o���9�Q%S�@��~ai� ���X�h��L#ܬ��l�$��ec�[ �\�&�v���ƭ,�߸�C�a�e����-�����aS'�4᧰]@�&۠ �L�R�=�̋� ����ŗy���֮���CbG2۾���9�Q"^K���C��j���Ee�6���n���DjԴWi���EV@��z�h*P���9��e�`v��y�R�8�a "Z�a��r�fŎ��lI{f��Z�m,���V`�Ӟ�\ w������|̗�l-�N~Vu����#;	v�����������Ƌ(��]Dٯ湯�H ��	��42q楁��������3��˂��h�����1��T��u��
0_���	���P�Ab
[�{��^ݻpmB2_�o�7w9
+�%/a%17�پ��-ۃcq�8}6j��O�r��Q�k�Y"r8��bn'}�q��\�M̿��|�sH����y�{hq�0�$�RC�����<��^\r�c��ejsAz��Q��g���'���'���b4r�R�K��b	ݲ��H�G��{��(i2ו���Z>ݐ�jҌ�VC�����R����=��;6�
)���Ɯ
$#K�� �9Ed���^�od��£�\��Α�?]�0vt�Q�H3y�{|zu�E�Ӹ��i�Z��yȵ��==3t�%���S�c��(��X�I�|f������u��p*9�r++�	+KOi?P ��dG���4�����S7��0���1�ꑚ�������٨��ur���p����S�,2���gt	&3��s���7��n�V�1�ELRmVԄ1��������ڳ.��K7�<1����0�7�Q��+<�q� h-!*j��壎h������h��k��S8��	��q���t���LS���ާ�K�����p7��2�����Ս�)���R�eT��;ߨP�����]Z���#ڋ	��v^�seI!$��37Y�-ɼs��b/�V Ay��"��>[猍o�B
9x]�v�����¸V�S�b�3���e:��$B�ǂ�ұu�V�O.65�-M��&�����l�כ:Ln�a��f�8^BM���Z��:�	97���i{Á!di�F
ke�؜�E��CG#O7bo��q�˥L~dj�g���?�	��45�A�B�y 3;��]uxs��!�=a��ܗÔ@���m��EK=BY̫����}+cr+��#S����N&�J��:~��l��An�,�[(���d>k?�_�Q��6�8izN�_��l�C�������L�0g?P}s]��P�C;������϶��S(�L��62K�(o�\���n�r�Ʃ�w(�}Wgg� Z��%�p�
ƥ��[�䶊��������Hf	t#*.�&�ayc�쭻�x[r�z7p�UQI̟W�v)dG�a���ϯ���C���y��Xb�#��S�R�z�8x"\�Z(�3{��\F��B��Y8�dG���.��̍�t�n�Wz|��Y��w��/��zc�nƟK�H{���]����abݭB6��zFf:,C��	l�?`���9�m���ʨiYd��8Rî.B���h��8m6�ӱ9�@��,�#���t�.U'�4��R�N�ᖩ~�(,�q��ㄪv��r���Ę�;#��]���0���Ҫ ^�ل��f���>b��� Q��Cp�L�����xp���5 ���;4��gq��EʾUД.���n6�c�����V�ԇ�= h嚔؆YN��P�K'�����b\v��,6���N�WV$یm�w�����(}�n�����
��r�bL%z�	�D��݂?,���	DWnGz��}��L c$\=�5%«��s�Z���-"�J�l�� c�1�>hai�:~�)���aݽ�T C�ȃ4��\��]U�,����M�,�
k+���>�iRɧ�Z���o��6_7Zq�$d�yy�s���fYL�<+�����W�iLM�ʥ:�q.���-�\������2���ͮА��BFG�|	Z����mᘕ["a�;��2��P��
ޔz�i���CS�&�Ƣc2�^�~N@5b��iQE���>f0�w흀��zC�1�D�R�6\<Xd����N���eb�b下�[ l����3���I��c��j�V8"XF���=Qb�w��)ﬧN̻�6��d�&�Չ"�T��������;�ҟ<E���b|�q�����[Y��^L�\�S��}��TܯN��l	��PK���4�ThO�:6�I���I��9R� ��l������Qf���#�:,�uaP�|Go�:xj�]0Fa`�Qtƶ~V���	%�Ϊ��Y����q7�͂hL�Mج���Oʐ'���H�pB%\���j�2�-e(��l>��:�`[��̬{y�n�ӼD�@��VB��~s�%���Y��R�\n	��������1�Jn@2�:��L /����NQC�	Zf�9u�.��`�����&`��Yw[�k�r��kiŲ]p�t�SW(�}�,a�hz���N�/c.B~�-��
C԰��K2�a
�	�� �"h�8'4����ߐ��x�� ,�s�ۄ�>��lF��A����{HX}�|Z��s�E�_P�0�O
X;r_-Q\�O�C#X묄�|�;���<q5ʳ^�V�k�N�Y�JR��cy"'o\"��"Q����*ǌVp�8���G{Lr�Q;�����>�Zx@�
�^���?��5�i����)��M/֧��RQo|>4��7����v)��I����Ԡ��t[��o������+�b �����y���G�.�\�f��͛-%�W�NP�?Z^����8,9<�*��y����������LW<g&qmz%��)5"�	�ȡ-�ԭ4�5.xc`x�S���FU��%��3���XG���uɐ0n�X9*�Z�?����e�|���k�U�gK�lG7���� ���S��j>�O���-��|�
��y�5[s~�?ыǴ��t�,��m��#,8u����1_F��n7QZ��?���}��k���6-��0��\!�WM�f�Q�SC@�l��l}���˧1�G~�Zε��������[��[OC�+���b���8�� *�1��ᇀ�=��nW&K�	9�06�,®�<���UBL2�ܵ�\�z~%��(`�N��H��&n�"(��C)i����}�9��Q�6�]G$����,��]�)Ϭ˭7aAwYx -�{C�h��G
!�mk�;�w�#S[�@D־ge�"���$���JV@õ�vNa�|��h�!�@��ԭΐtyrO�*��}������̏��yEmu�hS�fg8yӲ�,���dDѲe���E�H�	�Y$�l٭d*wR�Y��@�X�]�����h�Ƽ�;��х�������6P ����7&ܚ'����,97�@�CK��R�,6���w���4�ܽ��ܒ��/M��8�x�n�G�t�p�����Gsln=�n��s�1c�P)�f�~��K\�כ�\�H!b����(�j��(I�4���po5����!<z������
��_&���G�z]�����	�kbe��T�����6�P v��ɣ_����я&��A���hzK�h��[��
�m�����	�8C��x�'=��L�~A��<��Ȫ�a>���V�&v�*�"�݋F4Jfw�v�X^�Vb���f�Im}J�q[����mpa���3ߗ`O��x��$*�7D��Ϗ�:]y9�4�`<��D�T��r�S��x.�kuݔC�ET�l���=<~��,�NB��y��������t�:# W�yLR�����C�'�`?�[Qx�i�e�>�u������i��cBM5ZÖO6"0D��~4]u�3- �ʪS>�Mg"����v3̔� ��1ꞹryņ8|)7����3j,R�̺{n1�l���z�����Z"Mʼ�=��#��|�{�P�?����vI�b{7C_�f�V{���7���lC��rMOp��ٹ����o��	<RL_m��
����6\�W'� ��t��#�XJ�
���#�~�D�!i�^rՋ�����$5z���	|���}R�?
���;��Q��G�h� 60U$0�R]*���.���ך��sNt,��nW���=Qc���)+�z4�]�b���+eT��t�Z֚&x��m�ݑ�f�R,J�z�
U��C�bi0�
n�94��\��0]M��s6V�8��-&޹�-Q�5p�\�ֶ��>c���&�t�M6t�7=U ����<v�^����V�Qtu��\�.�^������8����1qy��d#=6<s�w	x�C�1XJ#(R�q�\&���͒"=	_��m�h�F����6��+��a�(w*#�zA��
�DXJ��pg�ZM�����ߥ�ˢhؤ-���q���3 $��
���DyE܀�o@�3N*W]H��_��ШX*3�I���(S�N��~�*��-j���Y��Զ޷N+䵍H�BH1Ph��l�|!:�g��+�\F����&�x�0}�=��g4����ѫ?�w�	Uv7ޅWp��V�
, CN��97?��qRw�ŨǞ.M�~�f��P�޲ɬ}��{��r�`�(�ILp������U�� ��;)�����墚�u�;���	!`g�0���
������� ��i��T*�B�|4�Φ�x��ȳ��N١���R�8к��^?\��mđB�����q��׎G���9�z2�`S2��bk����H��z�aJ��k"���fE#��R�̏�Hmf� n����̝��W<c.�V �˓� T��&A�C�P��Q{�����)E��L�/-���R�c�b�zs�O�eנpk�~�\#j7�iLa��l��i~q�LH,SoU+���L��7�
�v?�	o�b����g<�n,,�5e�s�`C#�8��rn��#�6��|�?�2�=*�Ϻ���M��a(i�ج��J4'!�[���>�cq
b���{�v�'^����\��T��2��w�M���ْ�1��|�V�>�>쏒(��u�/NF���f�bA3b�QW����ɗq��C��2�Q����s�P��������P1y7�:��R�kĖn;V(�`�+4�̛�%��mP�.�\5X9���ѥc�)�ί��1�����
������� {����x�;!�ڴ�dѾ��.��Z d(��o����{k�;~5m�y�Gv��E#�������8���T�k�%�h���Jg�O����g�)e �kY�$
v"��;th���x0�xY	$�s��g���S�OKD;t�^�VyĞ�^�3��DW�j\F�L����i�Yc	�@��=9�,G���<� z:/�au8���Q���=-5�0kV}��#B�K�`�9�Ts�%�͗fmk��s��S]���#���r�Ҥ����@�h��r^�ϭ�����A�$��A��7&acTg�74��%�6���y=C�o;�K�>Z�U�3��Jk�yb�od�|���MA��u��>tR�U��x\�;���u�8Y�9r�z��9�^jX�pV֎�3��9�_��|(���g��Ij�wdA� �����?�k�A��*vq븴��O2��������Pdm�:]�.Q�-��ּ^���O���S#����e�"�pK�l�r� ��K�W��A�w�Z5[�	���	�� L�%�.�h+�� ��'4w��Qi*8�9h��پ�fB���66o��5z9<�S�s�)�!��t/�#p������0��V�AbS�mq���=���g6O��b����s&?�4	1�~D���� "�C��U��(Y6Ӻi�~�9��u�K��싙���H���Ɏ��ټX�����-]�A;>�zBj�p]Qz�����wO���V���e�8,���rױ�ãQ)���ְn���[>����Q�\5�<R�$1�s�6m&���}Wi��yЯ,Gmv����%K��ñ�:Aȼs��y��u�-�h��]�C�3�W���޽��S� �.��BG�>>���ٮ��3�1�r?��H���̐@y�Q�������-��g�#S>_]\�Q:��v0�0��Zp�p8T��e��#��J����t&��,}���ܼ�,�k�
xu�N=����$j��.D3����qe���@l#�=%�/M�	�;>���m�}�D������l����S)��̴�����r_��#�D̮�����7��_T��j"Ք�=��
fOa^o�xEs�˗_׬4x%.�]�*G���o��+%
:#�E��Sd�Dg�x����۾���6���o���2��R���,x��S�2>���j '}��GU���������˴�����w�/j:��K&(���Æ�́-]�LB���5�7��l�^�6@�i���p��ۺ`s�p��&����2�0nߎ�Lv�&Q�l����v;B�ᓙ^�h�G�]��(�����R��P�K�=�N^��-b�/�1`� �����)���VR��.O������;XZv2K�x�h_��%2^����Ub�_�0�����X�~5%,\q�PN��P�S�|CY��w<Cտ#rhS���*P,jb@v�b*>��ܖr;[y���BFbZT��S_�PT��G=����x�e�T�͘�SH�~�~���_ꚒȥY&��o�d����Q��K�ݶ�2S9�>���	�]:jQ�4X^=t�xG,A��if�I��f[�i��\h��h�����DM"�tQu�m�㧯yHI8Q1�hU����K������0M�P�r� ^���"���0�J�xz���h�)t�w�X�3���6D2�6$��R�ݐGq՘��@8:�Az����i��m�w;����(�/��}�v��=�5���݄d�lF�����rz���&�:L�e�/�>Qb��fps�d&���3��ҙ`�Q ƶ5���E@��	zܣS$�
YEs �+r���	!�|�������� (G�f�M��)vn��w�	�]�t�ء���4�~o���/�ši�.&{A��� ���7=6%Di[�?�3?��dY�W쇌�@��1țb�}"�yY���+��><cё����?'B/��+�m�7#��������S���j�5�D@:A��5��[5I'�[�����vLE-��<������D�%"V�����,�^��̩J���KB�h��g�*W9�$ q�h��+Z/�˴�e��sH�j1exS�b�m7���c�������XU0 q���n���ݰ�ԝ)���'4Ƹ9\g��R�.3�Ӟn&QI��=�Q]ƅ��vA�����<,�k��<��#Y���� '#Y�9�=]�,�F�x�x^�!�.M	���#T�{.�F����rZ[�A �QmMd�{:����(��@\.��8�]nw�B�hz��c�*�[��+���u�U,݆�/���uF�F5��nǝ����[<�]=Ǎ�H>9\�����A�r�arHy17��jU}੩V��*�M�]�b媂��W&�iFO�Z����SI��w5�El����E#w��ߥ��(Q�J�?����Hi�	A�(3�5�c_-BJ|��Mw�n�.L��N�C��=��S�.��,>�C8�<~��7;7��j�=� ���*vV�,�]�j=��-L���N��oV�����Q�X�E�D���x�fdÓ�l��4��I�y��T1��Ug�&JK$�Q\��Ӎn�]�}��Ϧb솗�u9)��<�?y��`]�yR[Q���L}雹�S|'˰��b�2^o��~�5!�ډ�)`���8����G�M�����-�|�jX�^��:b����c����D�b���s>���+NW~�R�ٷ�O���z�d,�	�Q���O���Պ����m�{G��F����]$9F������R���QU���&�й�8�O)��w�H)HcTQc�b)��w�s�Rt�2uܑ](ġ`����X���v�L��>�'i�=i|te��n�����2 K����I�}�f@�d�G^�w��SB�QH�Zty	ޖ��<��VD?k��;Z����4u�� 0�9�,�� {ol. Bj���X�:k'�G������GK�	�8ɨ���zT���8KF��&�X��+��<���j� ֿ���:� k�������6;�4S�/�˴�'����[�iСG��'�6L�/��O/. 9z	ح�#Y?ף�n��B��� 6�a3�e
�v!#�դs�628&�8�#_:���ֻ�Vty�0�T:W�P� Us����>5�ШX��s��J�D����=��T�"�jsl�3���!/'�6��*%|�I�,oW��(y����ghׅ��#Z~:Hk�q�'���7�����+ @o�� �Y-�X��P�8������d�ą�{3���c�X�j���v>��%�9�{uD԰�:���`����uo3 ^gf�0Q�朖G&GN�j�|I���Mv�M�'�m�~�п�j40���������{Vܜ �P�_��<���-�ի��a8E�ix,���Ԭhƙ��jʖ�<t���EWr}��gU�k���C�nB�b^:��PQn ��`�����2��-���72�gR:���cx6��t`K�A�k����lyc�@�o��e��.������˻�A�?���vF|3p����Dئ8I]��XC�A�����o�uս�� �Zhp�[^k�_�I�i�������@2��N��u&9L�ta�C/&��������I�NQ�ia�u������_AH��b�:v �K+wJ��ݬj"g�\A>ii��.���VEk]�Iޓ詂��YUK��5yj����%�k�|!q���!�:�����y��j�|8��J��p���O[�c�i�ݥ]%����i�[Y�{7��9L��"��!���c"�e���T�^�Ԋ�ʛ	Vm�C�����p��A�a�4l��Ⱥ���]���~l���(�-�Y峒Փ�4_E@��9��A��/�.�>T̷�)�K�����w�u��_l5�ȋ��\5���r�|��,kT��!���?{ę�-�� D�^�g��qBw�9�RԕWq؄А%���.���}�#�X��{r�5��ސ���"�l�?VO�A��&�oP�<T��ne5 l���/�>��w�u��Jh�@Ud
�iHe-�������|��@����X������-�n�3�I�!IP؜_08��&MBb�W�c���^ޏ��Dn!��נ��$E� �)��Y��!-�㥽z?6�H�mЅ��3�����Lm+Mշ9�H�e�=�{���jY/E��p�"WjwRiq�AoO��=l1��n�6�c�K��=�}:B�@�ո^����94�C����ϙ��00����Q�B����
���peV�g��ʰb
b�2_OQ��Y��-�Vt������ʓ��Dmw@�K4���+��Ӄ;�$˃�wbu�v�N��iwq�P`x`��F��l�ic�O2'�.
�8vͩοg=<(|Nߨ�h}(��_�(����3R��q�s���y3��(�\L�%kԱ�Վ�Ɲ����	�Q �y�u��%JqK2R4[�\^�!��_�iJ����}����@7?m�>��eM3��R&���2�8-Y����e&����!�q���&�r}��� ۢy�0E�id	K��>A�+�dN�Y�ek�s�VD��5[�($Q�ĩ%b���Sq�:4.�d��ҙ��`�ai�~2Y8��
<��h��p�I0�����&W�%,5�����U_属�W�SA�Qߎ����;tT��㨺�G?�(�Cv ����d5ԤpC9��KK�-j�h�"[6Fn��j�L����K���'Z `S����.& W�>H�}5�0��U߷�rn�t�OH��_je=��-g��ʳ�(��>md���?_n�^�VZ���۹�vVPgbWɋ��i�m��,s��]�zv��x����;-������A�Ί>.�i.I�Ó�r��GB@����92��TD*�L�,�A��
]�U�c~0<n܏c��=������	n��}A�2�EwH�4�b����I��������(����bX�%J�6���8���"׶P�5��������T;Xxa��A�D�i���Zج���§| Z[6��S]p�h����k��W*�t�v?��E����5��`�+yx� ���wYwu˺>��ۼ'$��gY9��@�#�k5]�0��2��,�!M��̽x�_tq��G����15kfrN2�_c���³�S�c�M�h�¡ŗ%��wQu�p�l�b��|��y"Aks�4r-�0���(�c-��B���X����G��ښ3�&��|B��6E������.�^՚�ʓ�����*��w��e,��8��/��c���,|�T���݇��C�5Ϊ�1��V..q�]�<�WS-Z:���{�\ߡLrGN�a��Ź��E{}�����A+;L]��=����Mfb�Z��ݞ�+��F�r�LN7CBb�����p�A 6Kw^!���|�95����}~��:;J[K��	��o��8���C��5J#��x�uo�s^��!�=�����`�@ߖC������0el<�4d�4:�����G�+<"o�M(ϐ��F�鮧����;��0�e�b��qM�r��X2n'��!�x]�߫S������cz�=�����mC1�����IN�k���ykOt;j ,~J4�48XYN'�tS����Ξ+ϩ��{��4ұ�FtW���1摤U}HE�3�M�gCN����,#M�2$Y��c�T:�嶞~զ���U�L����
ޣ4���>`��j���f�|���F�׻�-l~�=ܳ7<ċ���pZV�<�(,%#��Aֿ̾���mCN�o{0�������D���<�çП������)ؒ�nd�s�B����AaW��~��>+�bG�%ԗ���k��a��o���ti$Y�≻��\P�M1��������!V�FS�_/����%�k֒�k{m����;�6w�#�����D��2bp��� v7���/֌��ԑ'L�r)�o����Jy���w�!�r��W�c���J^�lҸg\�cy���u�7�C��-npA
��$�=�&&d���d-vx�N��%���*��� ]R�T���/���|�Vi���{s��A�.6�$���X�]-P�K��E)���WiwiV�Zݟ���/�����؉�P>�I�w�<��od�4�z����$E�ÐbF����efH��o���ci����v&�)�-c�o�UE6F�8\_ڍ�o~z�w5��� ����,L�Z�q�* h��r�EL��� �`P%J�[<�;b�

&�ѽ��~p��b�>�"Д��h���7E�]���I�d	�>A�E���N� �z-Y���s�Vd��o��&?�N��{���ܲa&= ���_!�[Q໒E�\�Y�x���kK/`���o���5~��%	�j U�џ
ZU y[{�Z?��I�4�&��8y����8c��nh�i�Wc�vrbE���h�s��nQ������3�:����i����!�����/Nh�?��A
}ph>:H���t����N�Q��T4��cD��yR��Z:�T�8Ls[*�Ző���KIL�@�T�z>�Z�Q�02V�!��r�5�R&�',��xqF�%���Z?��g��]�Ї��s=za3�w�םώM��4G��͏�2�ӣ��6~�i����t�Kl�z݊����ҩ�$d�<����J���*�WC�4�"~�"�"=��|�5	ϛј~��P��=,���'���{���[K�L:��uJ ��it�F�tD�`�)��-��c�6xG�e��X�[�S�K����x������&{D�e0��Ym'M5Ԃ�a�K���^N�[2�5����B�4y&�ZI]�u�\N�o r���H}�׋�9pZgg*n�T;�-�p�;FJ>
�U��Y3�IDr��������8�U�� (o�>�5x8����-5S�y�m���^���h�����)�=C�_�&v,�1�(H��\�Q*�V$F�l1�
�ًb�:��k<$1�b/��:
���/��@dM�p)�L����}����QCOW��,�
J35��~/J�٫+p��g��s�����.�h^Hl�8R�C�X^;�~��ne��WH�f�6�X�nR'���g$[(e�1Fu���9�c	���H��0jNY�/������(�}����[ٶo�R�샠�3�S љǀ}fv)�Ǥ+�����"���!8�O<���
.�Ӽz�H�.��yOjs�� �#(@P9l(�v�����˵����MW�N�^ayϙE�K���=|�~�< �i� �}&�3	�z��@5'��`�oiat0V�]����yTݩ�a�~�����f�����"/]���.��*��U�朽k�П��{f&a�J"�*��?K��=h0i�s��W&㔞2�*{��w;V�Ҁ?��7(k���u��Z���R��o�e��j2��2�Q�o�N���. 5|#N\�J�ʷ�Y������U�_�6�@<�}���VjO#�i���۩B��0�Σ�7D�={��Ӫ�����0�)��eP�{���j�!&f6,�����O	�����yq�.��
��GtMj���K�m��1DS|�����QC7(��� �hi��!��]4:E<z��t��'��wl?!/vz��~�K���/�H6���aY$8��a�c�rd��#�v���q�&FWo3��ky�d���_��������s�s�Q$n*�4
Y_69�}�)���`��$���|l�(�Y�îDL�&�Cp����k��m}���\���z����/�r&zC-�_��)��1�<�8�O>��Hbu� ��������g�3��Q�L���깟�aI���{�9p�w�'�k�ewe��կ��\}��@�]�Nv��E�L4j�e_#ܶ���W`1`h��1JK�i3�@��U:�FO|Ux�>�
>ȑ���(<9������)���-=f��꼀��u?^�	l�P��[���ߤrL��z��:���&��L�Que��Q�]O�n(�&��+m�]�ޟ`Xq�U�Z"H#�5��d��w�!|�^	�'�ͱ�Mc��B�