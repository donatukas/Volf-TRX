// DEBUG.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module DEBUG (
		input  wire [23:0] probe  // probes.probe
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("DBG1"),
		.probe_width             (24),
		.source_width            (0),
		.enable_metastability    ("NO")
	) in_system_sources_probes_0 (
		.probe (probe)  // probes.probe
	);

endmodule
