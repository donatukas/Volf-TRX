��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.��Q�"Gx��F���C9y����.��@��l��omCF|>7��-�+��z�q=��y�	�`!B��J��b�"�_?Ʃ>,���w�f	��ħL��	�Գ�]α�������>��fܞ�T�ޭ� �V�,/�R���eϡ��ʆ�m44�O�r�{hj�D��KH�J�(06�ݭC�O�Fd�uq���	ad���u�hN꬇����a��+蹌\{�%���L�P�o�����MPbf��N���K�:�nQ����9���.� �έ���sU�|�]S�B��>3c�����_ԯ�=�<��{�^vԠ��T�g_kф���)��7��j-��G�}��[H�}����w�s�9�9��+cL��&`�m)^3��?��y�^��pKa��=_����	(�O6���I�C�Av�A� �v1��7�������2;��h�`��`��?����K�P��D����gv�k8nS3�C��2ms�A�bNe욨�DL����,���x_���
�����!�)�����A�J��ux���m�Ue���]i�1%ըA��<�y���8�z�!ұv�b�p��+K9�RǾ8����|n8Â�z�pŶ̬�A�P~�Ұ�c��#���,��Y���oP����I4u8��w"<W{R��Jfb�k)i13�Q.��m��:���!�$����o}�8'�!���e�'�����k[M	����lE(�
x��d��w�`
��sh܄nj�����������*�Z5(�߸o���n<����=�N�"��lV ���x@�P&�w	 ?n�T\�pR�.\ �б�:��1H$,+�E�����Q�s�}�1YR[���_Pr-(X"ע$x�>�����{��BcqX��������Vk0��,O��'�Z0���NmE��p��a�tQ�(!7' ��0A�ʳ��i��4�<�<ne�^�����
0n��}�ԅ_�L��Ƹ��Z/�}-��o\%�{�Tb�m��/�¾�n5c�zOt���۟E��6/��f�`�����j/��Z���s����z���:n��;�2�;p��$��p9���o0I^�h�%Bv��)���l%焥�ӱ+�fH}�g���'?�D}�a[y*?�Z Ǧk'����ɸ~Ft�0�z��C�SR�g�������隯V�b�do���m������-���%��[;�;ͱ!&�*:��ow�j|�v�9'XϨ����ҏ�@�n(�`_��<U���s&g��g"�xՒMQ����~�q4؊�g���;ɷ8�*W�>�x&W43���!�acgY���8���5Y��+�#��'65[�m�uR"
T��u?�l���nY#�=繜ѿN��o��L�����0C��΋$�.��� y�ïoIg�|{� ���ȯ6 ���B~���^����x�M-����{���yTs7}�&��^B���|Ep����0tO|"�C�{�m���fs�����;��g��fc"{(dH���1Ƙ�u�v��0����RS�����GHr��1�V�BP��kZmN�%� Y��zh����Z�F>;7�����9O�5by���峂L� ҃$�2�	����J�a8 ���;ɳ%Q�����՝w\�D4~U�g5ҷkԣ/H�K8����E���,k0��`|����w������v9�L�̭��}	�("'떆zpV��0O��dNi�������0�HS�஗Q��j�:l��H��]w�$|E����׺c�e�moft2c#��[^�e8Q,`��|e�^G m%HHe%Ӧ��,E4!���ًE�ٱHQ?��;A\d�C�[��f�x]1�ڈc�И�o���{������x((ם�_�����{��0\b�:�d������ ��&��,"��*s���qOxJ&���w�U��'��Hn�p��~lO���:��e��aQU���n��)�*��)��d�� �:�m�Wګ`�T+���YF���cb��c'h40~/>e�7��^�~`4V�
Kq?�����.F��N�-'\�f���fU���I�c��R����{婴��3YI���'�r�k`�g���	�҉�>�^H