��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~�f�?|�ў.mh� M_�>/��zTg��P��Y�@��+����t����m"�Q�e���VW=I��K�'�n]�	5���	a>PZ�I¥��Ԑ0���^��r�s��)uD��>˯tp˲O9�U�%���h�#$�Ɯ���Ua��+��cO�p<[�������`=�eH;y��,K�]�#b>�6���Y�з����M �%�R��P��dC��}��(��ܐD$�_��
S-�wM�_!߅l��Ұ���k��~승�,öJ`k��r�x}�+����/�>�� 1�KP�L���}t!�Tğ�:0�/�|�ry�eKQ�l��CEv��L,2#�t���A����4�(�~g�a^+�'��"�9��Nŵ�D�̜3v{�|�*:���nf�~��	{[h�kw��=�
�l���KIq��nT��#c��t���pu��6Ǹ����:���.�\)��t�V�2Q��z���^JL11�����ɠd���m��b�$��wt�K�Gwq�t!{9�)�v�H�3m�w_�)NӲA7�X!��xu��LR"fcOߨ����x���n�AV@+?��;�L���ѓ�s�:�5
VT�p�U��@�'A{��V2H���F�|Z>Y�K��K�?�)f�0M<�����K�����xW�p��R����2�� I��tF�B.Ĕ�%�֢�<s�E�V���f��Me^�E$4�X07yqG���'y/{?0}K`8��5��C�������*�Xp�v>,<H<ʟ�(i�d)��;�����T(��qN��!Z3�ŷd�>@�SJ����S��0]0~C0>H����K��!%�c`���ß4i�)�1�>�z�'_��/ݻ��3��V#�(Y���yEg��׌�	�Jl�6��v���1 ͫ(ix�kvߗ��Z٠���W�B��[�����-� ���rXO�`�ȈH�Mtc�
��\]����z��u�B�
��7�
����.1�*�혗�s�q���6EڿK�iH��+�58�Q]����ޞ `�ќ�����Q�L� `|B����ω�����y��.l�n8v�0ψ�¼^ꦗo��L���~�M�K�����V/�>��+h��"���}��3�a (iT��fN{h�{?��f`��.��nBUg�/���9�L����� &��b� �%��x;y��l���v4����D�����_7����,������l/w�y�!p��0Ҥ� �I�)	c2b��@p�����	�%iF��-8�>}ۡ�eRΏ�1�S��� "+��C��FD� �"[�~�j������fҶ&ʒ�<bS�|Y�)�a�K$����ٿ/��",��������6�7���3l/�1Yaf7�s����� 椉�����9��h� 9��s�<�]����4�c��kF����y]��	b/�_XNǕ�}�}�ֳ8�`�<�ª9`#��yg�>��X�x�J�W���$��pp�{c��)�SAK���x�%��t���vYq)�e?wn��ſ媛ӆ�ߌ� $��R��8���d�M�0r#�*_7m"���lZ1���iqX[1���;�$4�gL�3�ζf��|-z�и�K׬eZ�ܙ�[�O���0��+w&���@3���{�,Pf�� k�������T�(A����J�xi��=�����؍ac컙 9����]	(鬞��9��rMպS^Ѹ�M�)�͏K�}�sݟ)<ڐcYrn�	<
��,��<�j���������%�D#�&��/�x!IdO��o��=𿂍f3�1g@ƓX�A�Y|b�r��{+p`$�u�L!J]޾w���K�P4��g�H[
��R���׾�e������Z�p�-��A������*.U����pm����9A,�zն������P[�&�AS��i����A;��i�������uiI,�T���|7'�������f���S�������A<*P[ ���G9�F��3��Ț��t�!�plh�
$�{�_"vI�c'03;w�>������H�M5��V���LF�3n�T�F��8��9��S�H�H��1ѳ�(n�h �}��W���{FG�Py�����1��j�_��j�a�w3���"`!���su`B����������q�w��#��d�!�j	f�ܼHOiH~�&�������3���9�N��s��p{��s�^{a���D���==����M��(��/�[#'2H?�El��?E8f�k��)$
���k���;+F����.�������\�Z�9��-�y*J�x���X�6	R^�%eRލ60��Vl�gR��i�����,���.�Q[��ʖ3�,����.Ʃ���ߛ5���}��"��w�I_V#�4�NgDxLq$RBŁХJ���~��&�H��Ipb����]��B���@L������7y��*旼��\#�O��Gj�ɌZKMЏ,0T��6v�y�f�A*S��˯f�7�Y�f����~ZZ�[����g���!��C��0v�f�H;�,?�����4���y�/%t�
X�ӡ�cຫi�M�4bP3����|����Q�lb��P��o:�0���y۠JU�_���d���|B���pRm��ZO��a�8�5��2����G���g�7m�1og�X�L5S�yQ���1�5��݁Kj6>���T��	��m�s^�2\Y����ą�&-�G��	����� �gw��
J�5Yc6w6�+��\>��F�@(�V������O��Jfd�ٝ]�I�|u���Bf���d��-\_C&Ԋ���8X$$XXӟS�<����e�a�F$�q3������q���5����XoN�h޾dc�f9�46y�A^����A�QhÑ>�-��	��}17������	�������G����K��
�AY+C;��ޥ���"upt�to,c��h������s(x��58P> 􄓮��w����,����XCo�ez�,Wez�$tʥ��QCQg2���˦u"@��#ut#gX�²( ���5��F{��z����[^�J���Q5�;u��!�{�f�{ï���t�_�g��n�sO^�zJ_nQQ����l{�)�Z�K��QucL�w���9�.�8�z����Fc;��v�/��j�E���l�:%�#���x�w��}A!�O��T"$]^������#N
�ǲ�Hs=Mev��FHqb����#2"�[���� ���WNar��q\w+
� �S}i�l���D��#M"+M=W [�,nRΜ�QY
�-M���й(9��B���2����fNY���N+�(:y3sv�B�Gh�*��Cd��6A�vG�W���4�*9,
KG�2O��^���� &������R�:1�R�h�H�N�\��븹r�p�6v��L�����Tt�mR�@X�8��2�C�V���y��h-�8ICgxj�R�^
����(��أ*ޤ-��o���j8�R�am��w�h��"�R��K�	.�7�ng�Yt�d��⽮M�"��������S,<���,kmW4I!o�F9Wf�B��.P� �k��^m�X�#5v')?DW�G�؂�lJP�]�lǕ CK���ΎVr�:2�a����I���ο�t���}W�_S��w/��eE^���!އ���@,��_���#��P��W���\m҃�l|��N�< ��9����I�������@6ѧ��G���b���8g���@sE+���/�@qŴo�U�_�.�n`Aޖ���%�f��Y�V�B����ͅ�ϕx`�r ��Ry7	�>�˟ 饮��I��ec��樮�t��@���Y�4ُ�J���CK������<��m>�Ԓ`��ȮSL��N�M��]oD�ņ�W.��d����vȑj�������c!����5�50v��t�NH���Ģ�[v0��� �$�� ����=���裟���B����u���J����4:w~۪�u�J(�	�n��O��Лg�1$�S��,�=T��{Q\��c1���0��d]��̢u���%r��_P?~�}٧��d_���&��:�GތK�F�����-Ъ��[��R��C�؁`1]���XCxx�����w\���ؤ��_���_F�#��
ʉ,;��>*ݯ_�i!���#�;���_��k��w/�
_��|K�7�`1���~2��P�5d�cf�����e������_���5���ǁׇ�_s{:9\�T��<��ْ]�V��ﮫm=Ә0{��k�Ż
�7#�R��f$bg���^�6�^>�/Џ���ߗ3���=P_��A�De��ɰ��N����U�$Aûoi�L�w��Ў~`��l���d�s^&�������-�ʚ�g�!n����i�%:>�������w���L�@sA�T]�]�T�H¹ՃK���l�/�J|�}12�ݖ�b��c�M���H9�ZH�)Hd6 Fk���5 �d�U��VN����a"�_ E�>����̕Q�&���b�^Ը��#T��5��BX����J`�l�~����D�ۥ����Z��c�$}t�	l�U���yA�9��x�*��4���N�5?Y�Ͼ��1�Y�+wi����;AX�seKu��ʥ%N�`����'@�r�������֋uw�a����\(��8�nȩq5��us��U�<NV�T���u~��	4�aP�^%1�'�9��
�*J��q�@���&�- ���vCTZ@S	�H�ܮ[e�j=��[kuJ�:�#�d3�l9;#�	��~L;r�D���u[��}$���1B��Ѿ9 8�i�\
w�b�^�'Wkf�n��3'���ɒ��3� b����K�5;i��ic���3Ͻ'�(�4�Ӳ�ʽH�:/�@abӼ�QJ�r���xޔ���:g�bJ�{�}��r`X����;�U��1l��h=��e6 �2<FU1�Y������Ck��6Q��i�x����	���!��K:���Ї�f����.i�v����pܹ#C����uŞ��/wv~'YE<�#�x�r��I�{.I, ��&#'f�e��CA���`�f��;=T��YH�/�*��x�?D�&�`IX��c��ީ�d��&�Kö��� �W,UsGx���:��9��78d���L!��$ð� 8����"�U������a۾M�ݏd$��$��}�;�_ߵ��$H��fD�a)��p~`S����~l}���5���`����ܥ��R�u<�~}VW�v��+�F�����E�˚͇{��ѭ��u`��f�@�bhC����%��{�6'��%F�Y��:o�bs@$2�[r3�S�ؐ
ؘUwכ(̝�Z�<�yF�	�Zh~�������[ �q|��x��>��dgplL�T���אq���`�X�k��C�n�T����/[Z9�q�,F��K����|R]Ji�7�S�o,�LN��l�dtn�ʪ�A�:��8"��}����n�Trs+6���U4g"�,�T�� �u`#a�<�p+������@@�](�����c�v5�z�+����C���bLu���D	�֘\�׽�&��wX�JR`��ϕ�t��w�52mo�q5�f�!	 ��w�?L������X+2'T5n�;� �G��	�=�Ri��[�B�|�+܀u��w̠�
�� �6����i��[2aχ�Ǖ�f���K�E�;�����_��$���"�h k�e��"F:7�>�Y�h�j��N���������B�CL7�+�O�dcx��2_�VL���r?�p���M��N5�h,~>E��YZB���儦��ۛ� 8��� D�=@H5��70�K��p���$*��ҀV�ka�P�`�j=�%�����p{���!	u�TK�	H�|���,p��<��&����{����O�v��T�~��o-X�z��&��y�O��Ҽ���%�U�Ky﵇��.�\LE�]IA��N���\�4���_��=��0x#�RLhN<�e�(��k���j���<��w�~�f��r/�/�� ��c�װ�*`�X��B^J����n�vc:�h�� ��t�oh@�'�=eF$�̩��x?�Ž�czK6n�)�v����B�k���)��W��P���_4	���c�4�1�_.�T8�I�W�{��j��x��rӄ���e-�"n��B��0�~�R