��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~�f�?|�ў.mh� M_�>/��zTg��P��Y�@��+����t����m"�Q�e���VW=I��K�']��GBI��|vz�ٸh��?8�2փ�%+.Ht���Ĝ婒e�])�5�Z��yRUn�M�����Y�?�8�>�R��2%��y�� �%����*2l�o$'6r�A[�q� ���1u�Fe���r����.�d��@L ���@��n�����Ax\��r��ق,^�h(�a���o�� �7���	峗�,�wL%��a)�?L�A�W�d#̜xW,�.#W�����K�"�d4,���lnd½��d��L̘�D9��)�Α�Zg�]��o?�
F�ؐ#n� 6�����\K��G��ܝ�w>{�:�O�<��e_�.I��a�����p���j��3�13�)�u�g�IW���x�-j�~ڤ�0yRG�����Db4^/��U+;�7VF(�M�.f���,,�.�$�"-E�?�RF�`ɭ�cYS��r�'8x`���ed��q�S�Q�h�oC�5Ʒ�d��-U��-ř*�d��fʱ��Ύyh{{���Ј-����-��r(�k�gn�ew&w��;G�0gY��H ���h��{������ 3����WE`dq�/����v��$��ʟ~�\���c8��L@߈p��ms�K�}x�ݎѫ^�O�Du�r�"Z��;�̵$� �1y�Jl�(C����!���m�!OڨR��D "�P�ui�
�*YXٌ�(�^�+@���$cL���	9��Q�D�3x��:�iFUW��������b�#Y�gA!h�U�����r@- ̵n�#*J��=6�'��f���
�[��{�E)1*���eR"�ٽ�]�`��Q�i�7���6�F�w���I�5�����+�R�Ν4������Ҵ�
׿0��#��z"gq���)��eO�fmr�у��yĠ
XY�T4Zk��WZ��-�8��{����Uw��f6��M���Vx��:$,��*!��+�aij_��� Ț�����@���^���9��20U����_k����a�_��q`潬F�X�vw���5�7D�q�<O��,��!t�h �O�q���X��F�� W��O����W��	m�.$�����@�_��b�3��� �y=��{�a2�������O��74�Y]A���\C=�tS�K�!ب��T+��f�e�9�Jյ�让�?s8�$(=�F�o���y\�Pj~&�\� Z�B�z�ʒ5��Z�K]5�~c:��[�����P��{������*�.����#�ɺNj�%�)�/r!r������m���	*��YH�~Qd��h��{�͹�ģ{�/ŏlr���,���_�d�m�U�i����;+q�ў�q[ ��H��U�Ay1/�Xo�L
.B!���h�E; ]�l�$#\d�B���q^��H��q&NcBV`����7���j��ӗ�L`�=�H5�����Q���S��ADp���b��6r���~�rJ�PB��ք��w*��Z�ӄ6�J��̯>��\����C��:"������Y�=
�	�崄G1<���b��6��ĭMN ���7��O��U��ʭ�#���EIR��PWo���@,a�:���:ph*Υ�gV�\]�c���h�5<Q�����,�`(9@�94�Vn,�z�=��z�u^ -��7�j+��^��|�o�C�)�.!U�%�Q�g�(;29{h(�B�,f�������y��Ϙ�E�\{!��3^�w~�HM���PS���SP��:���a��-�6-sI�܄:̑�8�®N�'�p�{�U�U�%.�C8<�6fj&O�.���}9G�s]0���.#A����2���4�[�R�G:��Ƞʴ �k�՝ә>0�yu�%e�\}�}Z�׮'�A'{��G�O�)��,�'[*U��wن��U�*Z�{�=l�/��Q�F��gb�\X�MvwI	3&���5� �272�"��<q�˖[�-o����c�`1˫����a�1����&�zC�[��2?�
���}��V<�����S�R���	�EZ%S��R$f�M�n]2h��$�0s��ǽ OdJ������A��\��T��������NuS;�I��G��1�������G��7��NN�*x�x��k� D|�r�)���C}K�,:�#a��ʱ��ˢ���jN�ne"��~2F҃��[�4	�$DuA+x�zh6����D�?j*�l/J|UxE
f�3��ljx�`��^�2�hˤ�!$I����p*9����bA�_!}�܅	u�A�i�����A�l^^���'���f!;�왺�^�ߎX4|�^	����b�!�d�۳�+�J�ہr�I.9B��Ω9�$z���f�̕u�Y�\�z�BW���BM��ן�~g!�;���Aۨy6�����8�{^s�M�X	��n�KI
{�-5�Sӿj��i��y��� 4���z1=�C_նϻ�>�'��5چ�%�4�#���]�gٗF�E<���i=P���4#am<ιg��O>a�nv���Q�Ї�X���:i揌���݃�$���FF�ou;���'��0C�kB��I�%����:'���F��{ q[��<#�k��wg�&���ٚd�&��B�c����%;��PW�m��ޯ�!t4i�{��>�&>`���O>Kb�P'�~ ��סh�\�N���;{SgiHȜ7ŅW�T���%mx���K�e�U�����L5*��T��H31���|����`�\���ŧQE�J�S����e.}A�b���4�;�;�!Uu��.�w�Y%&��u��d�4�k��0�v��q9��I�՘ב5]#r�6��kR���{��֢�Q��|^������z>yю��� �p/�N���a��D�9˒v��z6�;���x{ླྀ2D�N�0��$%�7Hz��UҒf\�'
��<���=���E�ps�G���:[=�˲�����3]��)��{���`���ZE�5��=��W�u�|I}4r�u�vcZC���ٕ���RC�(��r�j�jfG&�O`t�����[N������G;��]
J��v%� �mRjV����.%4{G��ʋ�@;ԞC��!��eCih�@�%��	���l�?U��]J��v�4�B����r��G2>��3�G.D�2]2���f:���7��qx��?,�^�5J��\ ��%iFk����"A�F��_�������d��|�^�������T��=W�LP̃%�Vߩ�ܕ�cӬk �uip��K��NT?�E�Ǘ���zuC�\�D������fj��Ѡ)\�_5��wq q���i�����(�^%��"Ց�./���\"�'Y\�/�"9���u(.�\�d�\���5�t��O��;�$ٹxm�	��`�H*��a�6Z�ե��`��s��K�?�H?�jzn�k�AȘ�AM"<�+��'�[�'^~qA_w!��
p���N1P8���4��z�A�Z����|)�%��;�������DcS��Wi�I+^e6~3�XzK{��������8�ԮI����*S�Ҵ���6��y�	�X��:��6`���C���Qz�q<����s[��,�V���~ԫs�3*�j���\L�j�b�d]H"��#k��f	��Ҙ���4���{�S#�����\[$���눃2u�v�V�.�_U�@��k��A+�u��i|��Wn��h�=����ܜ�Dr¾A��p���" ��1�Bzz����<kg'1R2E�!V&��J(���W[�(��>+��8��嚖��䫥)��|%T�z%�d�?����N��yz���T�sR�D}y�.Ɗ
�[/
�x^���'6X#�[�D��+�/�����aUQ������Ĺ��g�F�Gۇ>�@�L�:��.���!|dFA�o���oZ�6QT�p@�0���y!��ʪ.*���	��!	�ȡ����D���7�%~וMҠ����Zw�*˕�by	څK#Dr��5�i_�d�����?[@NK]g�p�~���������|Z=�EkN��u[���y�	�N��m���"�R�U�:w�B߄
��?T��X�Vӑ���@�?��1_	.���91�G�Y��$�����z�J¶��uq��@d���W��3����2^T#�*c݇���F���t�a-��F��o���뺫7�S�OM|�0JN'�Y�	���?Қ����u��r�����ޣ���B��S����ƫX��� $[LO-o��6�R�'o���al1F|$�X��d���p"���M�$񕤔���es�W��+���\$hJ�G���L̪Zzz���O�Y�y��5r�@(|�,V���2	�k�*z��<��.,eJ���L0x��Pc<�%rb�O� ��%6"~�Y��k��+.�':��a�����}�N̾�΀ ��]�`Ю��]��l�{��7�'iV0l�;a�Ӟs�����A�~%��]xR�^s�jJ�~��Qj.�7����޶|�D;�Rج�Y@!3b�7�L��2� j�y�愛`X',�F��${-{l�v�u�5?���K�gl#�&�ƍΖMtX3�oe��!5f9��A���Te�j��ĵ2�����aU��<A�n�ٽ�/����.4�08�}b������Y�P�zq7�á{Ȍ��Pǰ���5w��=�H���C��jB9:��^n��y�vpP����+[��.���������G�9o
4J��>=|`��o��fjt&n��cd�=���kD�L��r!Q`�g.W����/��'��(_�o����f���r�K�av�k�'w3�~1�;�2�9��}q��w�EZ��]pQM����]W���� �	:��j*�~
}�K���X�Ffh��O��ԯuM�I1��̓YZ�=��Iڊ�K�Y�;��Tt�Q��=F�v�[�_��:�U���x�OٔT��s}�}���+�3V�� ��X/E�A&L�������=�!-/����YRzY3�fҏEmOc�2�!f��R`g�࠴�*��t�T��P�裆.�&=�4/Ҵ�")S�oA�O�����W��(�X���1��]ީ����:�H���8���yە��&�����8�5v���������x���>�wf`_��������)��Fi�U<
.���4$��ᬈ����ɲtt�Tq�Y��#�fS��J&����F��!��<K�T�EɎ{,�P	IB��M�"��	n����0�;H�#�K����1�v�B�
NH��ޣb�^&�E�h�7�1X�����R�JڦE�h��?8k1O�.��B�:�k�'��[-�[YC�����j�ۥ%iV�L�	x�������톗cK�=��|�Q��<���3ϳ��ugq!}�9ٹ>t�#�Zvri��0���hs�R���tYj�( ���>�c���0n�{{�B��`*��CC�����5��s�Ԣ���}��LbW��k��\�'գ��������ฝ0@���@h�P�j���;'DJ�3Υb�8�����z�����؛�L��L���G�&p&9l!��d�K&� 0�g > ��Ǵ��`U	s6��
���`�% ?J\��E	������.��|�[1=����"�J�YL�!'��zbS�[�0y4Ju��G��Q�cnȗFm�nJ�{ۧ��
	��W�sQ��	��Ȟ�ͨ%Et6
h38ђ.�f��˙�J
��lf�
6��,�<m���?�vUl5�j���]>�(\�kG��3�ܐi�Y�P�^7��>�%�2#E2��s�Ơ���4v���b���5�hc<�Awe�H���8��>a�7yh�_�w���G_P�3y�]q�+#���k%��� ��P>aWo^@.���)����⤁�t����ey�v�5B��3h��UaE�K��RV�3�#<Z����!s��r�D�{���A6Z|�.�'����N�w�wsYX�N�9��3#�S�r��ec?@�ż����������:3����,�]ژ�0jCN�d䎈v}��;�ne����A����n���Y��Q�I�ig����'��3��fQ������<�m���]*㼈4A��Ϡ9��/�E{��a,��Ἴl��Z���{�2�9�����\`���N^M��DP�?7���D���^fp�޶���z�`5�ь����%}��"�P]`�J����� ����B`nGRi"��.T�Y(~�,�f6��s�qh��cg���b}aq>^��2��`dC�#�U7gM�Vd���*��s���Z3Ⅱ�wC����x���P���	݊m�$�tܦ�:�1�+v�7%)���G8?�ö~�ڜ5-8���Rc���;�5m��8�%X��!A(͆$*&�hԤ����$����Ǧ	'V��%~G�j�ĠZ�x4�KU��̥c��̈c:��BԊ�m-Ia㸴%���eQC�sy	��������h�_�.B"����N��?*���7*�p�'/�(��#�@��..Dn�a@a�#|�I�F�2���~" :�B�G����C��8�D2�o/�َi�4p�7Vdƭ�S���RV�$i9��~.���np��3˴ �INܣWwVS�_�N5����99���@m%�#a�S�<v
!���oR,�����2)�HZ�����V�;��9���FlN'�����}���r��J.�Ǭ�ߵ`�Lb�tN��������q����ɸ�͓p8����Gx?�g�7���t�n���ac�[Q�״&�ϧӽ� ����:���L�I�|G�l�<�,ʡV��
�g&^ŀ��H��Q^9�c��ο�C��~	�ao/�[<�،Ş�#�2����໸�y�T��9��u��<ۖ
)-S�3tμ����k4w�?�+���Q�7N�Y,���nC�r�?Ϡ��_\+�>$��I?�%䜳��+��Ǟ���96��1�Z��Bc�S�%	p �Q�� �˭��!�0'��7=���d2#�zlh'��vnF,���{=��¦*�	F�����Y�Φ�Cޘs1-y��� �u�נ�
3����ԗ�Z�ӗJm8	K���x�1~{�Π*�x��gq�>�Y����sm���Z��0"�u9���4^�~h�uϺ������cx�l�_J����t�A�f�5t�b`$���HS�J*�\l�mE��@�܏O�"A<��0�q5:�OF�d�%vJ�,Ҝ�T����rq��^���"H��$��5����&��xIU����qru:������X�Q�����JcR��=��� ���?���[w��uD�@��U0���:����uu
�^D	(闫%�r5D#��ѓ�5�+Q�:�9