��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.yu�=�6'��4��f�;�J�鰷:�ذ����?�R������Ԑ�r��ZJ��1�8c�č7n��MQ���������1������CZ���E���^��<�8��7����T.�nO0$�MP������m��ݪ��2��k`0nՁBD��bYWo�2C����v~/����P\��N�Ȭ��,R���rHx����b.�z��x��˴�C�ya*�gmӼ��q�L��>�Zb#\�R���|��M�_���W��9��2v�uv�R��q_�Hz�~�����XT���AE�`�A_l���$A���2󺛬H}���sѦ��T4�p�����L��*��Ӽ�|���7�Į�dU���J����#�_�d_ l `����󘖄>�#$�jH3AV*���+m�Z@X4���S� ��ØA��M�2rTB�Z�:E�������n}���2�f�s���c�4{\�$nfi�7h��a�����5􈋴�zGƢ2vLyT�Wg�Y��h>H��>��$�����b̔�wx��&���S~LlZBLҒ y�z�ؗ���p$t#���"����>�]QQ����ع[u�Bʄ�����*�XS�4���AיP�P'��4�s��j��.��\��r|��ڡ#�[w������'DX��.|��۹C� v��bl3�S����p1�pu�@ ��]����ɳ��X!��G��A�t�{�������a��y+�5]����̴�}[�|�~�i�i���шJ�d�d[�;��P��܏�M�`�Ӱ����B����ʏN/c��d�B8���h�V9���z�*�YS��@]VJ�ܩ���,�p�C;d!�+z5��D FLŨ���{Z!ET��`�P��nkȢ�ͮ+G
w�+O,�,�(�HU�w'�7��������Ujǋ��;��mr4���E� ��U.P�)��ҽN�jn��G�)��7+��;֨�����-����I���m���a��%�"��F��L��p�C(MwP�:����w�V���Β��"w�����8@I8Q�4���\vʤ�`k����>&��D�6ƎX��@ ]��d��4}�����/{7 6j��-�ٖ;�0\��$n��\�Ҩ�7��gU�Q��G��e}h�����Yc�l*��f̍Xbi^f.Ԛ)UOs�� f ��z�Z��.�V	�m����ݤ��,��'aͺ{�>����@錯��M�"�`J���Cd�wnb7��H��w�����a�	^	����>��u������G�9x�(�_��)$�{��ĺ >�4��L ��G9
r� ��������  �����A�,6	���rptO�b��߫�"En���d]xnG��Z���%�Ť|^P�H��������L@�b�1��#��׸�C��A��SO�0v�&���X�w[�����sX�[�Z8/<����8��pe�iê۲��:,��b�N���p�u���y�%>�sm����'�>0;��x�ϐ8W��*�x�"�{����7_�&�z�w��0��d�9�Z���/�<�$�d�W��U�˯@�Eu7	'X�:�t�8�?�WA�g\�Wrp�o\�l�lj�#���ܓg�*��gb��k���R	�ʄ�^w5��=N ���XڃR�1V�����<ż�kWԦ�P��ȃ�C��B�<����s��)���,��w��,�>�N�d'Q� �����+of\��������xniӾ�/�/~H���q]	uh�yKR�{�����v-��P�fF�A��ئb��VQ�;g���A�^J3	�"ۖ���y�p���D�ͼ�j�q��r���D�:޷�Å9����;�Jym|�[��ᶰ�2��>�:��(9��Y��/඙���p�^J�x���TR�J�1" �& P7�D�uy~a2C��u5yNo�(���G���x����r��8N��=�Ժ+�����;��D#���[�}��$6R>�'9���,���hcήm_����Xe���$A+;?iͬ�ģ�7� г!�:9�Y���1����;%3�3>��۴T��ȵ۲��h:�|԰m�)��Iit��9�ܤk�n^���$����@���-������ӴH�*��)�x� O��H���z�9!*<2�}�޷(c��6\!�::���%'j٩������J�&/&��gJ��H[`��6G�j3X �a�b����*����@^<-�ߞS�$����
��.L@~{�ChGYm�o�g���]$q°��js"����h�iZ��e]`P����ו�>@ˇՓ:i�/�L��s�b9Jr#�Ƨ=�/b�`�MA���=g$ϓ��A�� �h�6�c2��0�뾶SX�ܲ}: �f�I����GYB� ���[����Zz�����,-0�a7�}��Fv~��d�ɨa�mL���	��z�����u��N;eNz`�"�*�f�v�����w S�˒�B�͌7���z�����d�͔�I�=%e��|���?�O�狸�~F��M�W��+��:������/�uO�~O�X2M�t#�ʱ� ���ՙu��Y�&�=��?�M߼��c{	�O���?�y;#�>�tO��2�:`�8�،�w�;^F�*������B���֫�:�Ř��@����+�=[��N�E�Ȋ�zU�ӏ%~��40�.*Y�2F��fc(�~Grڤ�r�x�����gKq�KU/}l&2�9J��=k�ڽ����<��?�	�"�����ƅ̖ڣp��y�l�=��y�W�����p��c�Q�:ض@���Dv2C�t�]/_���o�sm��U���J�R���۞�,��Y��r�ܲf_ ���my'�����I�E�������a�&����ʔ*	9�Xn��8	�lo����9~��=:��_�	i�54�T����=�X��z�a�i�`o�����|��iG:Q<�/����X�/�:	���R��z���y�#U����*�{��B�8��_�z+�$d@��Hv>U�9_/1�/��{z���?%d����]g	Ap���@.�����nZ�i�Rh��>��]�MJ����ҟW17�����+�'Ko�6��g��W���T"�[e�Kd�c7ܯ֡:B��LՌ�ӫ���Qo��X���kR���!5l5��x��ù�̺��UU�֤�
����R��"�r����3]�="�
.Y���m���}��%�m�bg),��JZ9s��,��x24� Tm�PƖ@s���M�|���/8t,��ְ܊7Pz�/��2u|!�d��v���u.���nm�Ofhuw,i�e�`�2� D/��}�{�D�y~û �G�n����U|���JI$;���E���ﰅ9P��,�����b[r���L��)����W��Yn�+;v%�+Mob��_7�U�۽��⍶��ۨ���8M*�xB(����O��*ࠋ�V����+`�\N��V;����zZ�J��������z#k�&¼h���4�=��TbS�8��~L����#&�3�:���yE�ྨE�����YPӷ���g��_���qO�f���\{�����	+]�&��ɑ���S�X��1��\��.ƗG�e�+tm/70�6.��_��\��|��u�Pˇ����=��f�q~O����\��C��£$�) �|����f<��?R�%V��]#ʪ�hլ���c[)Әp.�����n�"w�U����-�ج+#l�{~�ƍS|.����P��k�D��Ў���MJ�����U`��e�v �-Զ�'���M�)�
�����������<��~*���Z�)Ɉav�h8˖!�'�kn���(pX:������;���?�7G_b�.���xT_��7� $�!��l6��W�dN=&� ��G-	�`�.olt<D7�x6&��}l`�*���ɠ��{z�O�R?�62�����#��K�sҋ���|�b�����H���A�7� �bK��F��8!�V��@-$��~>���ȢK����������~deSڴr/�ȏ���Eݞv"1hs�z _#��cǹs�{���jݝ�������u��E�޸t�#��Q������~�����-��HH\�J)��vp?�-�B"�0��6,6�_����O���T 'b�3M�y8��Ul�w.�ߩ%�B�0G(���6���L���݄'��������K�j�ȹ�;r��,���;&�b��`�7�8�M9���d������w�OR��uJ�������)�����\����5Ir��c�6�!*; }b��p3�4�*I<�O����9l��=PfC����v������%;wSfK��2�?����p��@����&������S-����ѸTe�<��G��EMtՊA��p$���'~�K�U��)���Y���36�� �ϔ��z!0�c&;\3�����胿�U6�#�*�;+�����7֗��(�T�<�u.���@�pN���vM�������>\�B��g��vf�п����ש���:�A�z	���+@����	 �|�s��1G?^T�u\�\�!��Q�����qQ��g� ��D�zu�*��t��T3�e�^X����[n�#�p9Hڇ� ��+��=�LQ�1%�Qdw�\"�ʚ ؙ�����|dYGY����fu��F g�C4X�XX56`Qc��8TJk5{���x��T���[pİ����y���0�t��J�i6�Ƌ:�8!���D��C��bL��MG�.�Z��E�.�.��q]�4H�H�G"�U��֦#��vjv{���AR�vf��:Rg��T���hZ�5�T�Ќ�����6QVl����������Ʌ��5�d<�>IQ֌���>�m���.��sdKbP<��)� L[��_�柔�Ǡ*�4��ӂ j��Bh��1�.1�^\��������R��:�#>�`Pkݣ产䰺��5	\ k��g��.��InV�l����l�O��	@���ֵ�����tA�3� �pמo+Y�h�/�jm?B���AT��`�%��čcF:�+B].� �@�sM.w���vԟ�)hys�O��'�P�,�B�=#���#||�W/��t��[C�p���� ��~<�k��4��p�c��K��-���8Poh}��S�t%�KY���j.�f�c�fGКJ��B�Q:��n��a��\����ÕeW��;�L��sG���^��`�&c �˥�.�C�_���m;�	�E�w��� Yq�� ����*?k�s	����as���&|%4Ĩ�̃i�ޕ��<!���šY���i�B����8��E{��ރ\��cvo"�D��
�K�W����_�R"�S>)�1t92��ٽ)���aӣ�8�Ϻ�
�M7ܡ22�>�/��w>��{Gw�ԆH�1��_�ۧ���Y�<gn�價�	�HVV��6mV�]:Ap�"�Z����z�7���D��X��0H>!-ٔ� A�N�1"�}d�#������ݣ�N7'���K asT\,��Y��p��g�W�7f]@�����P󆱈�;Q�a�<�.�.R����i�K���~�2t�V���Y�\V�,�gh*�6�$W)��ud�ڻ�aL_��弛i��B��yэ��	du�R��m�f-�P�U��á�*b9�-B����n�j�"�3VUzi�޸r8�=-����4^&��5��/��Gm+��q7ٙ����<sh\_�&�(�pG�@��#LY�'�T��+��71��C��t���A��5�� ���,��Aa�>�޷ݮG3��Y.�v�@ l�z2�� ���	0�]�j�Կ�L1��0U�-��T1����2$�'Ɍ�z��d!T�2��tv�g����T��j������[��mv	@�,����������u�w�%B��ɹ���|����@ĭ �c�u�� ��|~x���9t����ɸ��7��͊���WՓ���}�N��,�����su�5ƐWB�.&9� �M�b֖�y����M��!���Vɦ��2�q���n�yέQ���`�;hz�_jm�fc��84n�lDa������h��� `��������(��&�M=�|q2x$>`|�j��^�'W�Z�wŸ'�*�n%h�u�Q��f���܁��aB>$�J3"1�:��;~�>��'����q�+O��e!���g`��C��D�Z����y�C�u6�j�D�@u���g�T��qo�lb������THǚa�!��O�:|ԇ�X�x<H���X�V�&K�F	�!����Ȥ��f�:�G�l���-��ʧIܼ
��������	�l�.TS�v���b���ۥt<E/����	��<���Q������KY=�?�Z��X�������5���2�v't��]�0{�{^	�U4�����*��R����AϰM�h6w#���r�N��)_~�H�0�M$IE���*Jq�� �r��򧐁Ϟnrl'��;�� �� �:4����*�fJ\�QlAp�g'A������#��V�E(:��+�i��L� W��i��L�Ԧu��]���K����+Y�D�=jJi>����R�7u��b�ٝ���� p��ψZ֑����ڿnq�o��B��{Y,�t�䈷�usOsTOO���"	ܹ�P@ �����Q�/����Ug_4�n���Z�����_!�K���.)H��� o)#���@�<P�ߋ(0ȶ���+5��c�tl�-*��k@!�4��E��ʮ�mu�:�c!�#>�=�TͤB4���Huh�n�s
.�td�m�~��y�Q�)��Uf�cR8T�.��I�w�v��t��2a�f����嬸��5����������W]�r-%mǯYFb�]�P�9�y�6�g���k�{�4G���>S�3�b$r���W���]��=��*�W�,����x�n9��&j��x�?l��a�m��{�,
�)Aom・���b�����Qm0]����-�vW@`T�A�~K��P���P_�w�zb����ک�Q�jS���2.@��/6[�@WW�nY�>���1\�����my��"���[��^�x��[�'x��4��63�pG�,�ε8��f\��7���ԉb�^�p�_�;�O.�H��j�]"��C[�}J���ڨ:�͈J���5rZ��%��d�Q7x��n��}�"���&,���������K_�����Ot��q�˔R��e0��� @<\�ݟ���BS'��s���>w>b�=�U��Ѝ�7Ft%�����U�aܵ����eV�Ç��ź�S�'������{���q$M����F�Â�$_���`Ĵ/�e��N�6�h"␁�'��>��V������S��ltSI7���b��	ɋ�U�[E�����(�` �";yJ2X֣�3�Z���ߌ)�~�IO"��t�+1��K\ߪ�[��=��%��	ɒ������p�m���8:X�t6p���a�x6VŶ�8C�A����-qX7����5�k��{���I�pk/�j���\�|��	0h���h�85�6�+���v��(9���h������h�`���u��%+���!qE��Hv#��m�m<��g��)��5�M91zۂu��8p-��^_
�.����[��p�X���}�����n�Q@�PpT������a2߆�$yg���>-�4�-�}+��A�V�%aː�E¢�AsC��-6�*��Jf_n=/aEZq@S̴�o&�6��iN}�Fh�����!$t�S�'F���u��1���܇Jq��*���w���I��P��Q���