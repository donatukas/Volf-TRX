��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U�|�.@�-�d�qs�X�A���d~`�t����m^��&��w�~��Z��?�;�NK��b�T/�\��j�-o�3��'��)7j�������wi�/�<�����S�2"����"��㺔��t��~ڼ�]�/\GN�꿷��g �x��W33&�gT�*%�����z�K�W�T��+��@��/�\YKFz�H�bA�H�3�Pm��]���=VU���J�䈔�K�
���4����Ʋ����j6v8dK����UB���Zщ[�C�����ؾ2�v� �� ��
�{;s�b.�x ����RC��K�a�^�w�P�������f�6�.7�fr�t�2e�"���Y��/*W�i·ÿ��l��0������:��_��7>e��K�`8$+s�'��RSiFbPV_��˂�i��=�W4��gcg��)>�{��J�_6��'/)�0��IC���Z��D�����qpc*1@��������~8|vV4�=~T���<�,�Jc��Ǝ�5�K*�ml��c�-���zs*`�'j���y�D�z� �ֻb���R������Y^O�y��~ѱ�*}5���������[�#���"յ���|Aź"sD���`��X(�Z�(��;���l�\(2bwr�wQe8�FrdT~o�=���X����6�J�s)��$N���#Q(\e�
��-��i��#3��fxfn��=�ݝ���o��i��&L1�h�P���u�I��>D�."R�8���H���P?vb�Z5��+�m:/����^Hu�'6��r%��]�*蟹dcn"�Ċ|+չ�ݐ@�8Ol���Rbؔ>QO����Ko;��6��95~�uG+��b7��J�N����}���e���_�i/��t[�wJk�3�z�����_�l���f�ʆ��d�O�
,�V�>���)	5V�DS�a����O~x�������+�#GE��p�}J~�j���b}�׌4�ߡ)����p���^�5�:D��=����=�2
�i)R�ˏ��#4��f]3wd&A�����[g&�6�8k}���ϊ�?-���X8�g�Z�t��Z�y'����0�I� �[�x�@�.�?#��e�g����;vYE��$�;�?�	Qn��ڟ.h�3�)����J���3���4��3�4�ޮ��;���6��{�{��x��+��;�,.�5����.�����:��n�}��7*|�uLNk�c�"�ױx�8��{cӼ]������DTw�4��x�'>	�P��h���
J�>)Y���LF<ܱ�7�92��Ҟ�%�>n6�l�:�%͐z\-r1��ُ�������D����<j�M���1�|ICQp� �����r�[FA���R G�0�R:��S`��pȼ��9}<f���[9p����p��&���F�"c�*� "�R�*�1�)���
�zn1V�R��1pw��O�P+��uA$��W4Jav��ǈ�m�İ��jC�0L��.y��q $��_�{7�S�Od7��O`�l�C�J�q��-����[�
6����MY����1����ר』�}�F�'�th,h�y��O�S��(���&� Պ�G̎��Я���:B��B_	C<I凩�`s�O2x6I��K��H9$h�D�������Tn�U٣vX,|�\Q���H�{�"��B�+�����3Yk9]�0F>�b.mN�"��j����`�4lm����|z����I��[F������ݟ�I�D��?�I��_�1�&�`�:/�Vw8߹��q.���J��O�H��u@��Gc��l�ӝ�Y���=�О�G\q0���}�>��I��s��)$���@Q:�I��Zq�(�hf#�g����0H*�Q���K)j�i���E��Qڋr��8�/��Lư�	y�!`�qxdg0Z�;>hr�n��w��������q�WT���*�ج��g	PM�`����p\n�|\%���quRs/����{@"�<��{�F� S�S@��nt�`LJ;}a��T��T!���d'+cz3OF��>����*t��CD밌V�+�[ǭ���`�j���hj�D���d��ǎ�F���;�/��e�A+�5�X5|_���)
hu��J>OR2׋NH�JX���oS��=���-W#��&8��n�ϓ���B�1T��e1��:i�P\̃j5���@���av��7��J�i ,ߪwt���*^�hO��f%����\�vII��k�G�>��+ȉb����D��.K���&G�uH�v�;��
�̖ڵn�{L�t�썖��CF�>�X�n��)�t�h#��,Q�e4���i�*�(����%�&�vp`�T�7z�Z���[�LF���L�t_�?���5a�N��vJ@k�ؔC��a�_FK��m�Ň�߀���Dm����D��h�O�{�<7:�#�S��%���Q5��g{!��ň�CG+zx���5Н��M1Q!��?`v$x���p%��%O$�~�V���Ay� wP�;Sx`I�C��nz��.)d��jJ?��S����Y�F#�ԏX!��ςMǱ[�H���stz��e�g���$Zr|"@��H�����: �&(J�5"˘FG�d�2�쭯4ƌ����wSȨP�i�Q�.��52�`ܫ��r�z���F�hd_��h���Q�)� F�E���!�!��ۼ1�C'd8� 1;���m��VTSx�JKW�L��tIH;Q�\���V��9w,AZ��-��D]��&��]Dz;��j`sk�8L�M'/�J����>��W'1�����`�b	q0Y�EZ�3�ش�
�y�N�?{�T>����!:�B�֊�a��%����b��� ��r��J�/,Z�ṕ�~_�n��T
*��ΊW�A�q�š�ټ���Iqv3���s�H���wlH,�l���֖	�>��2xv#��Pg�����W��A�ԯ��b���՚�ѷ ��U��ֻ��h�.�����s��06��5��/ �yI��lN�A���7{��k�����O��k�4	m^����\���U�o��'�1�(��)���)��1)�Q���B��Cy��Y�A��+5ga���>H�ץM�X�+��҉�kn�E�+��]��ld�B���䊟�m�٘z�z��a'E)"�Ue�	�-����7c[\��ڢK>x���Us�ea��ڄS���I�p���V^Bb��Kڡyׅ�s;����
d��ֳ(�U�qf��IF� �����ԣ���p�S¡�].k�����בB��=
���J
�~th��F�=�'��Q3�m"��Z�p���XPx��~~�-�\��(������z�h@)�0w�\zb��m[���#x�	��~����Y.�>+��(�Ӆ��`���8n���l���&�z-�Ǌ��s�����,�G�@�s�� ����&J���m�;bȂ�h�9q�o9�6�u^�f��Q�]g�QF�fNV Z@5�S�<l��{yH�.vL����;��|~>%3�8i�g��J�,�w,K�|J���qo�"�u3_0:r{�zg�*b$��ы�X	<`�q�1nN��j���2�	;e�%��F��?������L3��R�Y�.�6	@��?����v����U�#�,��:t`�J�m;�Y�
_�՝�S�e6]خ�SHҡ�|(O����v� D"6��s#wzbQC��[��JǴ=�d�һ-�U�Zl`�P�G��%H�#�!��benń���Ak0R�H���a"�nx�6C�Z�d$�y�����΍�lN���G�s}@/�ێQ/e6n�K��kS�Rx�w��-�=��I�q�K&�0^�I&��ْ)1�G� ���"��gh�[���h�.�	Ū���m罢>-g�j�VE�˯�dd?�b��cc<��q�/J4Y����ُ$��Ef����ب+��"g/��a���+�� �;��G�tr�ȵ�Ӧ}�Iw�L��8��V�����&��RH��8R��Wk��%�̈����h���B�41��>�dv�;v����;R&��aM��srX��y-<�V��v��
j	��r����7����������e=UIs'���4���aAB�@�;5�F9-���B���ҷ	10=B�e�{�K�YYW*0�"�"/�j��i�G�s��:���-g6�	L�'���?TX��@�6���"P�3�֣���P1x[I��˦�G:�=�?��y�L87���^��X��7'��,�¤"�Z��v/#<LBъ[yH��
閼�Eq�τ��v�ҠS�O��c�cp�ZN]�#���}%a�9!�����~?�%V����H���ܑ�}��:�>�-�K��?us)��),����ma��:�kO��]� ��"����B$3{o����r/�Ԧ_�T�:���/�q��R�{z��}\`)������l���*�ɡ�b�s�����%�5��k�xl-0A|�tKWӘ�͈�`�%U%,�W;�,t�@Q/�A��g%o&D(\e}�#pV�ތLB�ë\�u����s�.1K\ZU�Ұ�`��(%	c�7�l���?M]�Ŋ�F���SjT� ��8��q��sV���ؽ
�,�J���]�$b�ӛm�"�����C,���S��Gm�=}5���"�S�C��Eld�����]��!}ihY�ަF�ڣ/���0�(�n�쳫-�O@"@�;�#����}f��a9yqL&gnQp-�Ͽ/��L;�h��>�N�2���S�R�c0m9K�c[i�!eJ0�P�(xH�S��Qz�M��N#��#�J���y#��<�]I����`@��wJ�����楺�b��B[ʧϲOo@�����4��l�nC��n1F�Wip���#anl!k��!��2�J�����4s	gK
HX�d�x�v�lL��)s��A��ZNQ�-��SkS�ĵ�wH|�+�]���r۞<�T���#&�
�8�N��Λ1�E;�o�#�u�@�*�3%��� ?cwwߜ~�f������������L���ЙK�	���?�E:����}q2�0��,ܼ��s�9^!�V2�'(�Б ���5����p�{�Z��{jz߀���R���c�O���tɗ�s���h���?�m�Y�H�]�w'��ܩ�u�"]�~�T3;::t�;Y�eFx`1�޵㧿��-f��ܸ�=���nK~bW��y�G{Ϟ=�;���P�p<:�o���x	°�$,�I1���Js��/��M�Y��Ńha�۴P��8�2�w����05aP�4&�0#�T��1;���ˏ���_��,��tC��8�J{XX*c��;���ϲ"�H���5��D*�7x�so{��E�g�>Z��_Ӯ�^}��r��l�/�Y���[lg�3X�?- �;�NE� ���r�^�`p����Oe+�vϕ�z �V g����{���`?���3�Ȟ��*��J��0Q��"�/���x��`o�p�PCJ�6����ԯ�jr��<�<��G����X֞�K-i�@�|'��M�6H&,�2�R���M�u?�悵�D�v�F���?%;�ϩ�4�Y��NEm�
BGq��q�@j	Z�W�V��A�Р�ک��_jM��?_�3m�ό[Ô��+�TcΦs4N!Y�3�V�7Ut��oS^��� wq�?#r��VE���X����ӽ�\�e@�֞��<��z=���/�w�q!;	@F5��5���[%�S%YD\zK�M?p^oߟ���I,��q�I`%�����^�C�0@ø�%�h����.��%���P�>6*��%��[����D�R���'*lbo��=b���KM������ulWٚ�z7��.�'5���h����\���5�㲱 ����q������Gّ^;��ʽ��&�JW��5a����Ha��(���=������|�J[B�$"e�=���Ur������?U�7�7{�\�"-=:�}�)q[8�j�~y��+3�ϑ��teQd��m��*�M�Y+OI���r��/��%�Z��+�	.(	�����U�Ikg����/��7�'BŜ� �(,���R����-Jcy��yt�m�6��|��t!xQ�H�EnM�A������ym������0%�1wڔ =�V��ɯx�)�{��?��*Q���ϰ�z�R8 <v)!�ₗ_?(��ލ!����n�~��z���Dcgesy@�,y��b"IB�x�ܖ���P=wDW\���K�=-��m��+�OKk�9����W��(B��"��K��d��I��W�v.q��~k���E�D	��Sh��� �/�=���/���]$^*���TL��WvIe�YF�F�x ��%�~e/���@:������[�dz�܊<��|R'M�@jɲ_F�O�{nI�	Qk��ZY����9��_�z���v��:(�*����.�:�Ż�b[/�7�t�0$ѵ���o��E�����!fo.�ݐ������U�~nX	y�#��#����unNȻ�!4�V��y�n����j��|JN�G��iy�G�|Z�tN�����Y�6�����l$���
q��<d����zL�l�Gd?D9�%�폭�mCC�r��F@���[2K��(I��V9m>$
B�����;/UJ)����