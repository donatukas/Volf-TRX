��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.yu�=�6	r��B��y��3�ˬo@�_b]/ͿBQV�_�|T�!c�Ǜ���Dف��<��+4�#�!ڙ;����ܨ[�w��9�je���6����K���1e'�*/I�O��t��� ���;F;��kIa��=I>ji�F����Q�c�-�;j�hIvmCI>��p�r��"����*u�����X�:����^��T�ң\t~�h|𖌓X���[�W��oV�{Ua�Ɨ�)"czC����Fl�2��-��Ѳ#lya�|m�z����#�E�2G񢶋rL�����i�a�u���z������Gt2'A5K"��t�7�p@a�h�qnpq������O�>"�������M�|������m��,�4Wk�,nܢ��Jx�
���1�S*�XS�]�͌p��d�\�`*�LmL�&�,�墙�zR������$�A�C6Y��ǜ�}ԭ����s
:blp��"�x,��5܂��u�MA?��ư����̝V�M^{A)4+D{uH�s� ��My^J��hZ<��`�
)�F ;�+<�SQ�23 )���3K��I�iRW;i�T�4�P�k�;Q1�}F-כ��1}�_-n�!�ВvY�:����e#n��w�s�N�Ox[�����Z�v1�}ҁF���]�Zt;g)]m�)�'��t����_T�"{~S�j+��b���Ls��6/8�]i�f�`�N�l��c��H �_����<R��oP���?�%!L�=s�&>��MϿ*:ĥ��Q?i?�
�����������M\�p�=���+�,�(����P��?+�?- 2jF�!w��Pμ���c3&)�?9�t6��U�a>�\���z'7+{�˓��^���~�Ina�9jc-�o�9�)W�S�\1mNgn7��T��>��R_�7hxbvY<t�ZxJu���[u�`z��u��Jȉf,#d�ZG
o�)�<��U�����[�!�ζ��#� ��^[�q��V96a�9���6�N�f�]gL�+��=�N//���tY_�̘�K'�cҀ�/��*b`�6Q=d1	.#U�a�t�>=r�]�t��q����-+�T[~��eI�\��|G�(��5��N8\���`�U$B���\/����0ݝ�<��	�m���@M䦍4�(!Ѓ�<O�F��Ccޟ�[�8�O�e�	��$�qkG�Md��A���*_F�Eקp���P�����5th�hf7(h|~��<*��<�o�F]SJ��'��-MIxj�{x���E��;A�wG`�S�Z�F3:�^"��Ys�T�b�}�h7�4�d ���8Ě꽂3J5>�Р�ء�u�A�1��a�D��S+)(��_]��	�ct�A!�"�i\͂:%�ܮ�3�n�m��S�s���nQ��-�-�2���o��ͧ���;��P()�O@E��7U�%R�0R�5�M���V�t��	�K3��}�< =v�~�#�,q����N�o����|��K��Y)��?ޗ��}EPV��[����u�P� v&d��o�/��7'�L�(�i{�{70���b�⤮�Y�ܪ9#��9��6�īP����)���y)^��u�K�BA/]f���m̭�G�		oS2N���U�{��%�u,Gm�	ӛs_tKDˀ�,M��m&�R��Yej#p��L�૊2j1z�)� jj$!�}�'����h����H��3���Z+�b�$cm"rumCJ/:q���:h��j5�p�8��(O������e� [_>�L���ro�9�*�Bg@D$�G��;��0����j	��,{
��
-x}�U`	:}@���I�A@�)��p:g�%��,�I�Ӝ`0��8�����8x�tc	 2�T�s�h05e�W%�t�,8��VX*�|ʰߋ5R��_�+�W�jՒ}�������Hd�@��qH�P��L���L��&oL@�v1I��3�c:��g����B����Q�<�@��M�h9mL��}���T�8ne�p��o�dG���jƮ��R�Vk�7�ƪ��a�`��L�~p���zς#����ɟ!�W��4}��_)�{3}���Z��$������{`��h��}oY����pƂ��ol�l%X�#���_�w8���`�S�e��3��Hv�W�I�!'������2Cl'�i� �zY��\��:��	�$4���!#�ic�^!_xC�`�"�@����<B����BP�u����[��^4�t���N�d�Ze Ug���¤�?��{ƕv�KC�@� �})T�Dr'"�ClLT������c��?��"�q�T©�O�vw�Ǝ��S:��uR��c`��3K�߭�����.�{�(�7z���l�C2�p�.J�{�I�-��N+�|(z��b>r�pSk�g[�����{LY��F�zxQ����e�t$�5+�fBD�v�����l����g�j��c�����g"!�"�5lC#����7j�2,=�2>+���y{E����Z�@~����x�쩺p+�����H��O����џ��^VQX�0|=�; �u&�{��inݻ~�+ �C�b\}��@����1).y�5�jҢ�IWV6j�Ɔ�˺B���c/v=<�-��ӹ3v�5���ja���y�g	�Mw�d��|Ub�`MV�/�p^��y���m�:����%F�	��K�j��^���h(���j�?m��\K$ h0�3LH����h�[�:H��5�ꅥV��my�6v�m�m���T�Fi�����Yv�s0=m�4v�[�G/'���2�:ܩO?S.?��0L��&?5�w{W�l_g������n%{��g{��굔�Gu~�Q�+�;�b[�L^]/�=C��b��o��J��8�q�V�7�-�D�Z�m�Qn�P6��Y�]�8�rY1[�u�N:r�z��9��a��P�^�{B�����+�b.��U��v�������K�x��eS���WF��J9��bK�lQ���M��Q@��8�Z���L��\`ЅS���2N=�b~���2�g�oClm}�t=���vĪ�e\�Ʌ8X(��O��a�&J�Pr���7?���cJ��z���F�ܶ��Wz"39U����������i�gl!3��F}�T�2����z���W��w��#��A�e��Oڰ
n�Zׁ���De�j��_	s+�
8�1�(|42H��	*��@� �C4�]
���-5���<%��Y#@�y���ka��4����� Ͳ`*W����2�9��;��'�fh@	�:(��wG��H��m0QRZH�v�-.' Y.�㿚D�/��Ҧo�]Ow�A���b��.ظ@���+)���$:]c����۽�F��=/� ֬u���1����9����T��cxR��_-8���������I���-����pL1��˧}m;#�п!mfG��RI�_*�y���N-O�q:�¨q<գ��:P�?��օ�{E�� }���'}ļ �xao�xU:�2�Z4�F�?���n�RMk�&'�� .�,�ʠpZҾ�E���0�a4����L-�>�S4V1�!*�p����L~���B,� lN�AR-3ި!�G����Gg&ٺxhDLj��/�m�_���4���;-N+�r�:e Ņ;tc�{m?o�B#TEb�-�N�#���.z�����XԈ$�L��͚���� ���v���Y����[����c��2QaEOM��8����7���7q\� <9&j��
H��
�ߍ�7j�ںS�6��**��L.�;uuZ�`4T'�$�X������i%�>�X���ZP>��.RJ���&w/Q�5��9 -j�����~?��k���t(e�@2�z�x��D?�W��	& Q!%,C����z�*w����ћhf�`���`���D�r�0i��:�yu�p94y�-��y��1hᆌ�$J#���i�Osj HMT����P�:��ټ���I��f���(&�a*�dX��wUf�	�k�U���1�N���S�GW��6�G�x�zu���uvk���|]�QF�Y �&���O��	j����u�q�x�tLB��d�.Jp������lqP�#��,ވ�z�v�[Q_�� 7�_����J�'z�N;c�i��\��趞L�Rvm]��p,\����W��Bj��a�®���f{�����dȜ���PR�j+R0ò�cQ�^�J�S��b��$��p����������[(\�	7Z�L�����[EX�b���oԼ.�BuɝK_�pG�R�V�Or�!dn�ޣ[��I����*���E��n���X��� �F����&0'78�ָpe��LI���G�9��is 3Yt�UĔ3p��`?�X��G��Xw{�ʆz���褾���-M���o�������>�~�p}�s����q,�W�eM�Ng��fM$�� ?�/DV_TE<ߤ�pN�ԑԖ�u�mb�dKgM��}�e�c(��%$��Ϋf2Л�9�
P(������tE\ |�y��q���TJ�u�yYG
�_�&�?�}�w6.��z��f/l;ܥ`�ԜH�ː@���|�<".�8��j�d`��U1CҦ��[�/	�4�ն��5>�|�3ClN�Gb��a7r�^X���8
��[�gg��ĉa��bWtm�o�?T������]�:U#��l�i�?Hm}�@��~߯𺡗��Ā.RT��7`��v������Px����bW�[3de��,��c��F��*�m^Q"�5���W̆�}
���6�\��vU���&-���`��#8�NG���<f�s��WE��@KCw�.��)��fRu��#�����3�il�g�t�~�pOx!׬��;�Z4i:W��N [�V�C�l�z��-�Μ)G��>�Um6�MF<��]�`���^��Ƣ`A��.K�J�C���0V,D� ���o���[�K8�]3�4�x�k�΋��J��ߘ{���*�oƣ?���,ǅFOb���� ��JU9;��#q� �O��6�_�QK�%_���X$ng�Tj]⵳�;pBb�����p~̈́��d���$:.Yfِ����o2g�����qN �������&=`y�I�uFS�V���bw�qlF���k��Ŗ�?�2�LNP3f����8��\�Z�~,�!j�4���,�M�M9c���WLcc'�j-1@}�̓��@)��!*����NO�u�m�]����*�׼"����z~T,�S,N`�V*���/��K�Jh��uj���E3=<�ƧN{u(tKcD�v�F��_��ן�a��bMQt��ϔ.\�ډ�(���0����+�+,���@��G�4�;9�K@��������= "������\W�&(eY����B����6��d���Q&V/;!�e'�'���-��|�o���d6��/BϞU[.�t���?�S�t�x�2E��'��D�]�3����� ���F~���S��d�6�Z�s0uYu�'l!Ӄ�_ݻ\���F�tm-̬jש���A���$�䪡��r��p�@�	a��=�6M[�O�����4� �&�)���8�A���X�'���r$~Z~2��<�-�<:+�"q��=2��)�ںe0~gBEW�e^9��>�m����j�T%��`�y�kj�{�V*��.V4d���\�kd���o��
0ՖQjv��%_�,��\���s�9��+��D:�<���'�������e���Xu:"�b�:"�j�)��u*�6����3kN�RS���[k��@K�B��olY^�I���F�[(����g~�@=kċ�a<L.df�w�o�,�!�:�~6/���`�Y�??Xes�0ᱎ�3A|gȧ�O�z�9J/Q��}�" ��dc�최�Y�}[�a	�{q�È9'.uf[�]�:�.9��V��{��d첄�����%���H�q�=S�m�[&��Ժ���F�Q\��B�o��0��	�:Ϭ��/I��Ohƌ�Ej�Ä�ޟ�7���=uH��NV�Zl��K�Ii��t���@g�S���c�!.��h!�R�y��I8��Uhd^�+؎K[�v��Qv3�o%p�0@\�
#A��q�׷��aL���B�q��VR����$�����g��~A�=Ӻt}��6������U/Q�2��y"y��@?�{�E|jr4��:���R:#q�y��w'Ī��i�맟���pj˟��A�~�����[����]��L���!�%m���F
 ��E��@�XHNZͨK�kѓ��h��I*׶��Rt�KȏW�c��86�����&� 	䋵%���+=�c-��ToZ�%� Մ�R��OI7�/!���q
���BH<����Q`��zF�����sR�}"�
$�|�/�������L�Q���/�f{d�K�qiX^�(�4NN�I��o6Wc��f����0�7��ɺ�&�q��$�����R8����Q, ��O�A�����a��eƃӏٳMWc+}%=SF!b;�D>��5�j�1�G���5g'؊������`���	���S=����u�)���8�p'���-m�`��}�'�.ad��qS6��w�,u���3�%:�e����O�l�M�Dg��5D�d{����#�X�����XA0*'٣��&j<W��i"��e�=��6>p��e�r&��7�� ��+�_)���N�;�&`�d�H��1�qy���T��1��zI$@Cn�����z@��^�H���i��_�� ��SzZ�)w��q���U�Y��y��{�%V�8�e�rX��<Z(a��1A����xw���1P�Gc(�T�PZ�7*k|��Cs!�4=�n��r�F�2�S69Qa��Rʮi^�����zV��u��/ɹ�♮p2/���=k��Q�w�؏��Q����>,�ug�͏���9iFf(���pb{�UFqO��	�_*�t�-ZV��-���̐+�K5�*/.��7��I����2��]����F�r��>avڲ�?�\���@
�Nkn��d� ׽� X��0�n�Tu(>�mԓJY�L�m����yU��dr����a�+�l,�9*e�ܐ[�J��dZ�� 5���kNBk�Sf�� ���}^�tA�fA��nd��BJ��ǵ`�p�)9
6I�o��3��w0�p���"�����IKG���K�V�J�ۡ���7���@k���g�gJZ�h�&�^�G�4��YAҩ/&�����"��+���*�{�� �~�잮��˖���<��.?�\�o�L�5}Nd.�h�nR��x�):��<�pIg*T�!WL��C���w@�o߻ge�ϐq�p4{�5h���� �/�&�^�>UAa+X��t��z�<T�@C��nx���8H|mN[�N�@�%X/$��D�}�0���2�����,h#!��de���Ψ7'.�1Ғ�pܵu���C�R��4|�+4�j�nF�ړ�����b(�HW��[�/ԅg��d���T��"�����08����D%蕍/�B;��ꍷ�u�]g)��f������ �Xþ}�X��>��q�R�M�9典�2g��P��;�1t`�{n���9���Xa�&�'�󉏔2lo�l�1 _��O����3u|֩�S�nP4�쮕�>���i�UxP������j9Q~�ު�0���/LA��'���AO+,����8��3OS�m��!�Aa�A<�P�z���_�&I����N��ό�C�Vx�C��Y����.��%���SO����6ˈ����&|Q�{�F`�v���&�Y�����OYl2����-JHp|	џj,S���wʥ�f�b�s4$�@��o�FXrW�\m��}�Ƞ�����N�u�f�~�ca�՞{<���\*@и	�����&*�(؆2.�F����� �k����+�����q.�;��E��B�e��Z^i�8b�m�4�Dc�9J�mn��1���)UV\yUi�X	5����� �;ÏJ�#�N�'N�ԯڗY�Zٳ2�]'��5r�)�?h�@���
K�D��JP�ph��?I'��"`�B�e�&��\����c�!�yO"��s"��找�����#�����	�'t(��{��rE7z��ӟ�C����Kߖ>%,����XM2��������a��GV⌉�T#Σ�	�~��6%��A�}�/���w�8a%��aƃ1��F�TRj�<x���U$���f��2�Y�ϔ�-���� X�����a͜୮!�?������Z
�$_)=��;��^a�J��˳I2t����/(^�vH�)���ci+�\����Q��+�✏��=�".�	�n���꘺v� +���6,����$%�T��sdt���<�Ȝ�lk��d����l���O��Ȩ��5���(����۝����V��oG�U	�׾մ�dU����0�{"b�|�q�৪��l���!��6�`���h�<������.��6�'� ��f��]W�-�9C�QfUAx�:V����;�iXB+�ݫ~k�{�t�1[%3uхHҖ��vN{���6'Z��\�(Q�?�� ����ڔ0���E�*�T�������e��8�.!���@�ix1���g>�c��lNd���+�&�PO��{}p�ez��`Ա�Vσ�j��$f�r�����h��3��݀�[V�a�͸�tÑ���F$<l4��hY_s�4\{U#������'p�=Ʒ]S<�Lz�6Ր®ʳ�[L��}�%�P��
4�r�（�=ţEzW�@��l��9�xDLѢ.��� Ѷq������j*y��^8ɿ�k#�E��PT�~��:�9��Y�7��d��깒�E�M��^�F��2 ^:@���Ϗ�Jk�t�-b��)��⿗�ˢy�U%���T��h������aͻmC�j�0�Z�&��#�Ums����͛Z��3��Y�p�D�k����3�vH߆�^�րA�p�tl�`�@�+��V_A��!R^û81W8�\�=�u ��H��S.��Sbn�Μ|�Q�S��@u���S���᷂���7�e�|w�&�e���bg��Q7�������n��1x�e�j�scP�S��fv��9s��OW���n���ܨ�{����y؋�y��N��W�WlR3��&9�{���G�K_��&�3<|���ovI�
c�+N�@����b��%2���9��8�c�Ҳ�Mvm��I��+�Rֲ���q�^����K��l�A}%�}i/Z�v�^�"�#�7���x��߼G�ʩ�E2q���(o
�y��NQ�@�09�B���	��ײ@L/D��~�o>Ʒ���N�|#;�5tԪ6�2�j��>	��&��3��83Y����R����-�^�O��R$�}nb8�A�Q�)T��Y�2T��i��؆���4+�ˢ~�33H�lרsyn4UN�Y�L�����AngI�:7[�+V�֚i̿�boq�f���.+TO�/{c�H��|& ��� w\?�\�n~��b4����AR"I�N:
��6�2���YIꪩ-Y���נT���:��\��h{�`}ğ/�~%$�(�삃B)�������ɠ�����Jխ�5������Tl&�vSo��[�U-�{CX��$�#&vh�S����teNQ�ol���^��M8�3¦��ygx���(D�P@e��Q��B��:�x�Ԯ<���z�hw=L!t����y�"A�|$� ��L*��߈v4v�#z�y���^��
u"Ҋ��{nW?��b'��G��s����y��@� c�@¼Q�j=fE���QwZ4r�	�ߺ��W��n��.�!��n�H��^���&�)K�`"��Y��h��d�����=b��M5~����iHM���Nq^Kqp0��_��W��&�i�頎7��.1R,7���`���������Vf핈0���XSL���Uz��9�26*J#5�����tX�0�!(G�	B�&�)�t�4�{�RՐ��?oj�fTۆ��?����n�Y���0jeU�0EPex[���U1.k|�hyb,�c��O���H�Pf���,E>.�<�_P���m��!��;��9����r8}%�p��ckpg�;���BW@�3�1�HՌ�*�w%�#��&>�׀�B�b�~׋��2�4���µ$��.��D�.����u�пCE�K~��r��	gF~2��t]]T#kI]�Q�}����Qp�&�a��V.�ݏ[=�޷�"��� բٺ�r���z5���J��zk��wla!��n1�D>Ҿ�#��6�ᖖ����/&2�/M�%H���x��6՛WB���}x�α�Q�|O�#�*k\J�*��뵋�ŋ61t2�vFU�q�� Kر��/��1�+x��~�Ҭʧ$��F��)M)�����_͏J�E�I-T�M�a\Y���H$���S#�&.���N���� Y��L8����*%�JEkq��6�LA�S�p�ᖰ�'��V����Dm��@��w���xP�6�y��b�
9������S�'1u����h��%S�T5����N�IG�����:��2���,8iH4O��PPi7��<�X�U�������6M��r�@�<�V�I2 �}����=q�rQ4���|Y���/Ł=M�/�͖`���4���ec|7^�4��!���y�Vap�Q�+HЧ�/�!Ӂ��s�,�[a�Y����QPT��K^ي¦�hDy�V.4o#�����_����e�l았׿x���+~�%�����TNb��k���� ��uܑ��uxF��`�4�u01��I�5ԟj�@8��t����X��7�,�%��ז�15�>��:a}0�Rg�뷏Q*t�xTWhL�)8�~��f�1Ʒ�y���2�䣁x��?�B=Χ�p˟J;أ��	/��������I	 6n;�m�+7��iw���s�sX(&O�U����Yn�����y�Z�P�ǔ�ˉO�>Y,-@໱ׯ`!u��Tަ��fޮ?;^]�A�ܾq�ͦ��o��'48�!�ɉ�" �+|��_��'V_MPL��Sw-� �l~/ݏ)2�)-����z\C�,�G��F�y�[����T��7:�P��ʻ	�?8a�b�����*'T(un�=��ƞ���g�%+�k��A�C� ��Tj^B��[޹'�|jVU�����L��?�D3�/�l��^���
�C���;~&eh����6-�ΧC9�,k��Pw�%�Q8�	�/-)���|�*S��Ԉ�����9�	b�h�ҕȒ�I�S1�R"3�{Q{v�j�`\��#07�H����F���*��p�e��@�G(/���vc��jƵ�G4��:唉c.2���!ֽ�������{�|���J�(ۓB'ٸi���&�(��~e��&�7vep4�7�<Na1�	���}��J�/vx�#u�� ���JI�i�ߍ_��$��)�F-���T��.	RrN�;L�»����p��1�����ɧ��ZvUIs����zn�^�>�����
�C�'#üL)[�x��q��~���vm��G��Й�=d@.���]�r�X
�9�M�P!�����Pӵ��n��U���UI��k�,ŇfT���[ȉ�3�I��J�d9������,���5d��N�R�b��H!�(���D�^vaȼVђ��V\bP4����U�����y��P�1�d'J����!K�q���`�G�}q���T(w9�^���Ny.@S��)�i�[�uE�fh�g���xv�6�Ȧ`?��H�L��FP0yrjJPf��WNw��O��}.�5c��:���5b�מt�:��	���CZVQ�±�2�O*��]��
��г6Cl�5��?��?�O��E��z]M.����ѓ#�J���,��u7�Ŏ! �[���4�<i7��{���*����>�zJ��]��|�*�hPY�W��K�S��,s�}V�'_���7נGof;DE��s��׫�/V $oY3]\��:B�G]�n��a8��Ah؝N���.�6���N:H�b����������ܔ��U���[�*B��R�;QMR,`�����LCOb*" e��I���ѕ*���R�n&�A<�.P�f�|M)6�6��"1�6���/O�R��"�o�N���\����ÀH��n������
i�����X�F?�fjukRU�=y�U��@��_������W��r�o*���$Ű�0:9�-#&�@�f%6���a�!���)��?�h,�(Lu\�lev��c���#X�M�rs� °�İ����bȐ�HX�7�@<%�@�Ei�`+���V^�.A��B&��_ݟ�zW�0|��!�H��E�)G� ��H��j&�����an��<ҝƸ!�3���+JMC�2�����7��<�^ѿ�G|�X,�ˠU��U=P��$�1��M�K��_Ƶ������B���z0 �"��F�DrU�0���>��K~u����А	$��/q�pc�BF�
�J���q��bT-2 &����%�^�:V�G��E_l�w�ʖ'�H�:H�ۏ�����S�~����m��=J#�%ဨ��dX�g�t^��$a�j�I�����B�8
a)�6�~O�A��7�8.B��c���݊�~���tl@WK�\Or���R-��U�s���(����[�s�J_�8%{C�5����t����eL6��z��en�jR^��4�'n���o5�`�.�����bgw����m��*ﲖ&���:�W�Q�H�������y �rl�uqs�:��q��D��9�2'd�@��q��H���l:�h)���+���������w�-�ӳxȋ�a+冢S���H��9�����NS���V��T��k��4�s6�w���6w���y �����q���V�z
���$V9>AX�gy|���;	k�����f~�(���� ;�h���	1J��b�H�A���B���<�{�{׿;��V������?��Џ�t+�``d^�d��[�+` �6�.%�|�57o%�=�`q�n/L�(;A���J;D�ߦz�Mq��^��Fe�(�D�DG0��W�:e	W�3��gU��ܬ�7gJ��� �sU��8,ݔ�R8�Oc�_91bߩ������=�
�d��Z�P��,�y߶�vc_�2����%?`�͎*1�.K��H��U�F/f�K����mג��;>�u2AE4�D�ϓ΂_]I����q�"��8% ���S�7.o�7�U���\�`���ܨf����L��T��{�W�׼C��#:�5\�_C�_�j{\��-�b�od'��y��"��AT����TJa�p���0D���<���a<R���Y��%�k6c�t�oM������?!������i���٘)`�D�2�y�_K���ٙ(r�Y��pP
D'����K�W�J�]ŒAPj���I�	k-�*=��� %~�Nx���e��A:�.�sB8#��Z>!h�Z��51U�&]��,�ɛ52��y�'ؤ��l�fFI�1�w#�ģ��*�֣��  �`x-g@U�He�X�еkSEo��P)r�Y2@HX�9��I�z|5#�B�WC߹i*��T���]"��R J����$�a��	��%h{��&�iSU�A0�	�b2�vn�k���X����Ɣ��C�0�a$cE���"U�2���m|�K

a�zT<�
Q�Y�D�i��*�6CU���e�_ˋ�!�c�`���u��N	�����Rfm]l�]��M�L2�ܙ=��zZ3ų�S1��a�0;0���MAۏ�lxr����v�Q��S�\,��Y�_��~&#?#�@lE�'֝f���ad`�}���'L;�ytח��ڣVX�(:��@ؼ�K���A�'���	�E&�\f��A�8��!h��;į]U>�א��>jx��U�y�pཎRd�b��H����Z)Ě��8�Z\����l��t��� ~�:k�H<�����BB�P��i*���j�����4ݬQVy�q�Z��&�~�	���
�g.1͑j��K%�ކ��n�;�f����"Xtp�K�;�3Bs�����H~��/1�O�-��r+ ��6����,��������`�hٔ���QA7z���(��f���s��eZ�5�� qC��^³"pFM����q���C~��S��vt�����	���7����,Bu�{��� ǈ�B�k�䯑�#�:�,Cʰqæ��e�n塧rj�v�ik���Ȑ�"Ъ<�A����A�2H�T�F��m`_|$"�8��r����ϥ�	߽�M��%\�-��wd|�pl�W�ܺ��g�;u�^������Ÿ-_y�k��1�:xU�j�x��b�S*�>��9��Z]?x��3���ԡ�h�e	������}{f�z1{GsC]��QsU��f�ʟ�5��ԁ�q�3��V�CR��1�2x=�/�E���3oN�)]ivu.��#@����{�H��{��xV�1���~zlgJ6s3F���Ļ���a���}j�	f�Ȉ��tA,D\���0���a�������-�>n��w1dyLS��L��{��R쟃��+G�%;G�*<5K�UXi���C{S��b�Gan"Q�g`�6����Q���T�_��gz��H}ɑ�j<�i68$!i]o�N}������'���#�9]��M6e?�D��Xg�?�w1�0�r�3W�\ �`��,��/Q\�w�Ld��N�ҽe���`�Fk+�*K��c��+�W�H;�o@�{�3����d)����� �����Q��Ҵ�e�����z�M%�^&�i"����}o��M1��B`�3M�V��k,�k�v|y;�#[/��`��wz�|����[�2�U�&N������GD�_K(����?�揣�$.�����9�����j�U�V��dN|�2���L�P�<�ȑy|�`�RH���Q#L��Ꮹ}�o��g^R*����1��hy�����h�ġЭ3�> Z�d�����),Js3>�r�?�
ZҒ�CH �՟13���*�U��1Y��i3��l�M��w]r�6�v���Š7�I{�����/ឃ?nSd��H�H����c+�yR	1�Q�^����!>J�Y�z��Il�(�5�C�"\B|0�/�)*��';T0sO�X��הK޽D��(B��h�"P&�B��x�0^�����_����}���!C��g�b��dC'��)Дgۡ�W�i�`[-P�@�Z�F�meM'M�'�AATN3�gnm�QԮ�y�h!������V��d�5%+�AA�<��1%��t\Fj�H�q{SA�C���'r�n�\�������d�fQmg���y��N �n0С�;��S�E2#f�'@�U��G�����#����f�N���.tb����~e9��Y�4a5�qǹ���#�ň=��D�%��g����r~��5=I�%z'�:k���-�y��1ث���œ�>������F!;BU0[޲�/��Y��ɥ�H~Ù���w�̖.�B^��u�Q+�49��|��㷎ϟ�%G��:^Z�Q+6�ۗ����~�]Ιl^�ʷ���A4{�O v������smτJ���/��1�6V)q� ��{�F�q����a�(�c,[�t�G����a�i;�k>���H�̧ǩ\8�����%���BOY�$L��Ֆ�\�i���.�9bU2�l~��DC"Ϟ4��AC���(�:���P5�����J�a-�҂z�;*��ydDr$�Z>�%f
�Z4�M�FCt5[��m�R�%��
�2�W��u����� 2n��)A�Dh��`����#|6 �;g�S6|�n��%yQJ�=�扩������-���Tp�d�&+�A�I�Ui��E�@ȢA�4C+��|�۠�(i��Rb�i�0&i�6H�U�2�!Ji%8�x$o_��t��CE�z|lMk�N��T�����Iw������ׂ��� br�":���H:��&uرN�����SӰ:��mW�z <ڬ����d/���aN�D��jxra��u��V�Ca$[4�m���M�s��}��'=�Q�#]�_���%��b���M�l�a����P���q�9�7���#�j��:8��OZ\�����SVS��N�5� 7؂��g�
�|h7�b����+]\�]�
2uy|1#���tNP�� �Qa����}�Sx���G�O����ez��c��M�i���@Y8�'�����<���u�%R2W�l8;8������I��y?R=D2A����;�xn�����C?���3ޖw6��>��:�GP�c�	-��׻$ߓ���I٧(T\����J��S�?����|(��n�tLaǺ#��qe�o>�-�;Q��J�,ψ��z��Ҧ�#�ݿb
��:C��:�hm���K����jO1����)����.pl^l�/d^�c�jOtO @)�g��'騨�4�6.�gq$砼c�N�?��M�cN&���x�?w�}�����RY}��X�ƛhגǃ�6i���F�]�iq���ї�V�+W��f�C��R���=�&y��D�[wy(�*���"���������p�@�@'u�������%sīٗ':�P��L/���|X��ػR��Q�k�+s0��H���gm���*���< C�I�.��tE獪����c�uưYl���u�9��x@<�y���P��f)A�1֏�O�w��AG�yߩ��B{%����(��S	�L���g��[7z��D����0n�`^W}��[mnl��U�B �H"�vG�֕�*�g��~�M&g�����$"&}QO�-)��;3\�����a =���1rp tdh�T��C�%P��`�=����>��"/b��H:s~�8�C� ɝaZNN��c]\�Ңp1a�,s�Xe�=ȡ6Y��p���#1�$*s�y���ma;��.x<>(����y+�s�_�+^<�IW"��H������|k�8���J:k,ڌ�C�����
�c���fN��Sdc?P')D$�$�ӛm��d�-��ij��o|c72��ɿ���3Ypy��3�/�-'.f��f>�A�zE��X���>�뇜 U�Q���o���v�i�:H��S�ax�Q�0NIr��g,5BE4hȀ߫Ф�&O�(Xs0��4}��V"�*԰�Q_NAL�A��F\�NU8��+"��;�\�*�b�`W��� ����^���R
�a�۰�9��r_�|��`��"�r#$��;E�bQ�>�ۀB���_脞I$���ӱ���h���U)w�B�4p�Y$�z%�������+EM: Q��V"}����5�|]��T�n,\Uj�Dy��s';
�22V(������Ƶ�@�6���Hd?9ȋ�[�б��1D��N2��(\~����[y��a�.7R��x�\�g!��yt�pS���0͵4e���"u������
�q�gk��姈�(�Q0��`�öQ0���:B����љ�S Mt /9���_W�k��оpH�v��wNSUԽw���W$���f�ǛE��f!�S;%�Tv�ŹB��[��dӊ7ԉ���08Մ<(�ϡ�f/�G�X���8Id�7��pS�U��j6s#��Hn��ic�u��:�ܴ�Q;��#gSN�n�2dI?2�2���������v|'bG4$���#�i�ZC'��^���@S�& -���˫��P}c�v)��W��a>����dp�Y&@OnZ�R�M���o1n�W
����7�a����� �^���� ��q��e'"��q�Z����G���l~��f��1�a8ts��e�nZ����L@��N�j
!b�ё��窭�U��x�?#$A��h�po��6 �L�X��
�+~?o���4u1��M\�66 �4{PöJ�ˣ�	��꧜h�ٟ��seႛ���U�)������ $s��i�:�4�וGͪ|��ߚ �����~�qY�d�ZGc+�2�6d�ީap�+M�Jm��-h�)��BL�}�����Ī�6<�r�.a���&���FV�Ipm�Fr(|Ĕ�,U���H��Vђ~�y�kޒM�R4��"�����ޏ
p�
� d�Ǔމq�V���ef�䆚��r�N5��e��fr�W၊��	;˧�4�'��͇���~�L�y{�A({�a���u"��w/��9��Z�IR�J~�6�R���=h��� .W�jc����T�g=��E�$���Ғ:�$~��1*���ƃ�ev��8잹�ȥB�~'��n����}oٔF�&V�ސZlR�jR�~|��楳&eR���#0_���V��bQ��>#�a��`{ڸ��/��+f m���%�����G�~[$T��\��=��l$?*lQ���%Y�l�i������i���ѡLꜗQlR_�v{*Ɩ֊w��p#d��bS������?�L�7�.�-�1O�RX�@��3N�?+N��[!Fw��&��-�2=�!qWnBY��
��u82�`I�]SK��0[��7#��s��o�7/�]�w6=SO-Pp �7�k�m�s��,�C�D����W��&�ȩ�w��M��hL�i򠌘����}�	�z���d��v�<%���b���Fu�N�i��mV�q�^�R��'�M2k�e�a�M`�U���gw���/Iz1#�b0�6�`�Ґ$��#���f9�A1�wsm#Uq�_=v���Px
���-�eO.s`&=�qDA^�E��\�\s��w��qJ��g'Gc{�������޵���0~�5�h`�CDda�`��d~,1v�Xiz�>H��m	��؎�D�B:����$�Ĥu�O<�*2�rC'� �$.�&�޽U�5M���S���r��J%�&7�O|�F�٤�{0_��'��h��f����z�+��k}󀧉��CM�G&�RXX�BuʈF�D�V�nu�w���������+
��͛�}��\��/�ѻ�Z��\��F��dw�@�����	���*[�k"i��7_{l�-jѽ��i�Puۊp�Uz+�9��GUgB�O�K.��q%��������r��ݯǇ�7̾p!��d�'e�;���ξ`	�$�3�h�6$�ꎌ�u6�z���eV�;���Al���� ��a8��: 
�b�R�AT�uc���'A	�K�>���Z�b��S��ŝ�E���(#���}}�OY���^���O�1`ޮ����Ք�r�~�'�zx��h��1;��+Z��v3v/�9�<g�HJ7_��X�J�o���=/u�lW�?