��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U�k�>�J�����0n�ߵ<$�h��.)��ND}��Nc��~\��J 4�������y�׬��K�8b�HD��[in4A&��ٕ+�Zx�d�*�w哣�N��eŕ�/��%n��q�)�>�/k[^��bbOV$�O���~�,L&vߦ��)e!� �41T�g��o��RG��b�(;�kPK%a)����̱�!C�W����"�\�y�'���Kʬ��{��r�٭�>M�.X	�b�Nf'dyYT�gWI�야�Hf��#��J����o��L5жw�1�n�3�8K��
��/ܼ m�]��%�+�9�΋j�c���o��]i<�4>����b������*��8LO�)y��� ӊ��[)x�ԧ��B��wM�㸮gK��I5f�zx���,�PB�h��c
��,ǫ}�����Ϲ�=U	��)���k��]~&�:~���w�_�j��u ��+�5J�V�p7�Y	荗V�%����K`��N�]�>AUV���J�2����S��O� ��6���d�A1_�B��a��ᖡ�Ӳ�$�و�0��1ƛ�DZ'V]��~�]q��aO� !G�Do:8���_��VHϝ{�t+;��-�:�}��F���T�����5�kH$l��k�B�\Uu���b���8M����2��)��#��ŚCˌך�Jmت1m���8u�DD,��6M�����W��6���>('�n���.w�#����+j���:޹���~L�6�"��#!);H��|�y�f"�s�A�	~�]����"�O�i(u�Q���-�:�
O�!�Оp��O�C�Z!�@m}�i&���a�.p0Z����:t��_T�$	��r6'�pZ8gǐ��'٧��ȹ��(~~�C��dZQF[�� ��O�Byi�M���{��4��04�������@�o�j��_�)l�K�"?l�&�s��S��'6%d聪C@75�Ԭ���]��3�C��*��"����r��I���D��Ҹ��Q,�H��@�ї	s_��ްi %�a_<R��(zFhd������bG��(/Ȗ�~%�N*���@o?�h�C���K)t�E�z�n,�ߴ΄"b<�,�s,�ْmR}]�k'��E���ƘO�_6��>�X�ٓ��T���+�q�9է�cV�3�_���f>q��r ?	=�L�S��\<���e�!�3�\w�'<Q'&��b3!�_7���"�J��#�o�$�����Vp����;>K�g���_C�� ��q/�� �4����@Q�}�n�9�y�x	��#���s�W�,�5�R.y��`���>Eu�q-�lA�=�����e(���Wi]�Pm�g�(��� O4�O��P/d�"7�D0� V���KI�Mͺ�~��v��q��Aղ%�L]a@w��>Q��7�ꃷY��t��e�jt�IRh�M9��XK�� {�
�]�$=!Su�3]A`JJ�xg>Rj�v��0Gm�6�c�3zU�i4�X?�7Ki`�
4�ͦ�:��6����Q����
7nj�R|�{nw�1hTC�B"�J�C��3�)�